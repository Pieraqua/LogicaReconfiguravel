`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
muhW37dPCIsOxWE/DM78T1WFPflrMc+jvcRURwxQ006Fj9S4ECJBxvIL/dc8YAaH
xwMc76bqlJJ7DN2uk+qyInnLSVkj7EpAtkSEkAhE+OwpQX5JvY8RjCYD3ZimgRa9
3Y+quSoAJusg0xg7mozuKeVaDt/ueB6xYlk9I2+sqOIHZsDu+CRvpNofTPPfkTP2
yyrlse13hyTG4BgRAs35gbfKivpXmj7tApIlQunofKA+Lju8TLlTQMgHISQ/9gOz
xH8alhuoBsTPdK00xPnrj0iJjpdvfNVhUxQt6Q+cLEZp84ePnyT0yvhUEa72AERd
8U7E1D9WuQ7loAU5P+Von8XLaQfEYQZ/9ttUgGQxYCNTnEiWr5JA3TKyPEI7pCxC
FLmtBDjeJxZbKYOMvMGtV+wqWARp0hPpmkh5fvAyizawLBGG1ZdDJB4YB20zX563
3vrrNji7UntVG0op6IW7TO+3HUma0x2rmoRWoHcFJCrtYN8Zd8GA3FlH/jQVFs/p
0ZZ+CvL3sgGNFEcCQ0saFdSlkoyXyuKIrmTSupAzbQ/S/Y7jRdNLJho4/bXK/53w
mhZFA6HlR7nO+HZ0nI+4jbCChTSR1K4HC449AdvyJOvYTVriFsrvEfR3mW+SdXL3
liXo1BcpeO8Ul7orn3G9KzDXkl4Ol/QubBR+q5T5hmIyTrCYndZxTYQlaljvjnEh
gLv3qkQQx1VNJ5OrfnG+ZHybCXPhytO3RqZqRXt0Y+PVg2qKRHvzKgJgqKtZTbcd
h4W5omAHB3sYi8NW3EGvh6TDDuJDUlbdkBjjAhAUt9uLEW++TmDgUI0jnRKjKMo0
dHw1V7u+4pWG8gds/ZDaGxhKZU2rKHSa2Yl9IcaEX5ua5BF2YC6ahaudq5Tm3j5K
rB9tX7saa0uaApxG83zSVYzB/tY6NACiXVXBR8V0XtbtKq2CgPGaDTsX1QspTnkJ
sSs4rx/XVP/yvkRSARwYDoBmk+S9u+NyY9/nB/LfPnsx5g2Ak2owHbuVD4dtO0/v
tO+mwyLN7FQtKdcHaia/0US19JEoz2qBIKZxtsMeDnZeZYpAVh65GXAKLFMQT+7p
OUP1rqALmGtO2OWL7m47cqYsjHP8navMYqDR+Xo7dzzMnyap7LnnLUSJPk43b5K9
Ny+pyLStra0YbxOeMMK2f0GiNcsBYnUEcQezvDAqaGzCkupfyjwslIf2nBsPL/rs
jY5rhFPuAkDpKfgD7VmzeeCfEcjrJcEhPtPnkqn7T/u9FAzaD3iVrh330pvy9raQ
id/mp3piiFHukQ6ucyw+XWcIdmO+ktuqOgbc5dvBIi2rtlMai5BUSUEZ9JlS1JQm
rYrXzwVqVYPEeOV6JUJ+mWAK8EnLGPofxU8TGV+Ocn+y2B+mIcPxikDcJvxC5jHw
B5nz4IC3emwCapgpzGXKvybOxcMCmERS2M6Aoqu5qy92UcffhrmMj65pdXCynckd
IG4wUiRUciQIjcpFJPacR/7MW48NqL3xBXZidz2dqJ/66qfkfWNhNmJ4WIblcq1R
8r8+Y91J2szbz75ii8jI8sL0mtijsrfAEV0QrjBh+up47yhOIoGBDg7dvVQCQ8Qg
R07mzPhttZ1RR4vgG3bHL2pZiuzh+fI4TATcD1+1VcFHlBJNrl1l+fLoOZYkG+lx
oe6ZZ4XWBgkENjMT2TTxxjrnC7kr5pHj0o5peQWgVmjmzsZb1TQfviBWjH4glOp8
+LywgwsSv5cak4ExpnY4zeCn5iV5VCsFhntoj4KCPyd0XI9crmC4vQHO2dcQQt38
lCtn+ujWpqLigXp5FX4AO/8u76Lg0+9iIdYbjsoY8SH69Y0cdLF/NNdxR5QP2nsw
WzgD4W/9qFUWBINgqn833Ex9mkoSmzRq47XjpKSLnl6NkgG1qa3R6WdvUOCUU6yB
qmQrWOEyQ1+f45uLLPwmBPl8IBx+g/+ZdSokxCq+21quRoEst2jHKNw1BB/5Ruhs
PSFvZwYPc8PhpBgaUyBeA9yQJQGP5D32sUlogpu1WzeG7m5DtQrb1elA9EhfiXnM
V4eK84mcVarNHXl19n3F/+HUS/6cd9eFU++mSbFw9s/d8J4sstBUV1lB+qE+2TZY
1ARvFmFYGHZDPg6FgwsnusCKgvn2iFwl6gRH7JRbGlyOPlfBbce141lwnduHETyB
DJqC2rqbS9xVK1hiaOxsaby34QUYA6w6beCFEFscQLy3U/nAFYjGyM2lfKDDH30M
jyNrSJpveDIgxywemThkjbntGvRugBcCg8IRf/UZapdPoFaMBcuFKG6ckLkejxYC
jq5vlVEtDJ6cG326OkJSpiD4DMJboGZqfiGTgTqYYRSxLWq5jAPp07jD8/ygWKYt
uGgVHD4VtOntL41uyJhjIDNGS3V2iaHMDh6mRJivPF98fCRGT8XJjvBNU+UO2Y1A
RUtRwneB2hAIWMq+oNNoyKk5Hi0diq71sW8a8GCKg9eYk8av9l6gMJsN+3RyWvKz
DqnAEtqotn1QUfBPrmAPylNA4gNqCr+zpsAXMvxj5kwkXJxqQ5foBrNtsfa3eoLD
7I4GigKcBPbqE6NgLkdQHds6OsNcz6I7QXQuJ2KCOIgKVXM5LmAs97Z5aP6ISKa/
CJjPsRqO8yL1XF/7/eXBDLKKpXYVZyXeDWon3ATs3oMFssoE0zd+tqFsJFSFn7J/
SwxTSwsPyhLyoPP4Ozd8iO2uMCVAYFA86xUfbYHDuJhya+EggC9bK1WY9ycUlLyB
KeFPk/CwGIca/3ivGLOSkeOaaMWDKIJEcaEO6w1gLRhq0rWej//FOUM26XGWU3NR
nd0Zod10/yic5+T2JclOxaEL+lGO/alzuXEkQvMPCjtHDUdshs0olOXlKi1Q2qQc
fHA9DUXpzvl9RkjgglsLavZrs+iFBy1GaKHESDvVVd6jdbbamEiKJFXXb3Wz+eCp
B4BUYG4kFCUAxp44g+JNBTRAQ/s/UUIcbF5Md6QT0MrI/hFRL6lx1rdsAIODZBCm
Br9gamJJvQom8k7wgxec5epsTzjLtW3nlQNAFD81Mi5PytzBnWmxDXV9KQWPHX1W
mmvQjG+nqzoEWS89i5lamU5tBwj413a+ra/czf7ZQt38jBORvMpiS4Cv9iXLrdx+
BGDzDczNw+oH+LTYitblb868GuliZPPHR0NfWNzExXJPf0qBI7mlQuDwkWa1TQGk
H4iFIwzUy5CJFjlTQlE2MPYpvDNdB7KyisCm8NKqdZil2ZjVJZbEfjO94VtT9EHk
/+s22bxm+tlQ6OKKFLhItrCfddrueqyytm1hhYvgx3y06Di207kN6PzQ2Xuj+W/H
tEIv1TPV+mBVAbAjiaBxGNuPTauybhVbr70xJwXrmUlu06vVhRTJ6GWoGCgB9mnr
eHWy5fi5zySQOG5ARg+k0NRgB/GIAFAojFByk+nnUdWRnp9RUarYWumRsbmub4kU
ErejTbQpzgApz2ngt0xCnMZUqJRVMk3fME9jOuYiUWx9Bx8+/X/5lsCtKIHsNAsH
7kd7w4NWJwGDiZ/AV9p/d7OJOlpzdMp2F7muoSEiWSGdHFebWTEM3yAcVuDEkdlH
+IVmkTHdIK9pZb8oBvYF19zZ5wvxjrc5z38UtGN3PdsN4R729sGn0TeKrZdtwjU6
YxqVmYqT1UprgJBnId5BFPvRLW0XhEafZEDb+qMfAX3ymJJlQFuAbkrNZIOzTOrx
3PUdYjIQlx9JVaUUOqiKdpMbsk2BZ9AH0M9os5HNsthfm/yfVx7gxTzgTpyVSGEF
H8waVupkeJG+0Odh+VtgqZnBW2eTDGQHTnVM9U7RVYqr6KnKLLhFggiJ3VRb13P9
5zHmfjJ6A1CFvnVlrboYDcMBU9VN+58OgaWEZ6US12X/3EcM7jL+XujtknDdHyvP
vkk9dVe3XwgA65stBqbjMPwbAOAmtvQaCNMX7EP4NnYNj0YDhXv9WBGLMcaAihng
wqJkQlVqbkogh4JS/doiGmMuJDcjnqC/rcHT9k3JtRN1FTy/lLAMUMNjvaUqzXnS
d4QE9mF2n/2Cd5B7rok9PmyKZ9n0Bs75SMe6d/fYIilobnNqb7vwTqADJrH2OSDP
8Q39pMcXmEnjyC7Ad1kNu+3xjmJpXsgn2nYUuXg5CP34CHQ9GgIzi5qW5Ifp+Hfr
9kC45k/uqDFYV9eZgsUWJ98sEFN4gHrusnFNWkUqlGgCSV1AK24VLBBJcftH2S+S
+tA0HE5IwFKXCZj01u5LGjW3/+hOEveQAgDkFEzdHwM/S2YTepHZAkj8MRdimeJX
IjL0LqiXLIGJ4rDLnyjvi7KfR8q9E5TswnxCbyhNiLXtbTZaH4ZECsYt6rNaIUHA
6H6Pp564LzUOiShvZW/l+HWABwAIq0Ocheb5RSS5Pk/ui6qyGz8rLIcqXTfZCQPr
v5pKHxJI3hAWOgOjHS1oLCU/I3Xely1t5JwP5fZzCgeTPFTv87/3A4XPD4MYeYIh
RlavKy8hN0lmws9n65Gcc5oYGajuh2ROWGEIeWioqzr91MJFCd7BtJjOHp0W1+NL
UJj2kywg/uhgbsAfzC1q3V1SSJtAJJ/1J9PxMwkPtHUvdRKkZ4O0TJqPpG+ReKkr
yTANSLC0hzYq6rRdw0Hf6b0hAG+AjfS/acG9tK+lwC817hRYTrmPn5u+R2znEr0y
ogGYCBwDCXG1/RxqrsdW6KQWvA+tF8CwCB/smTK9MfBV04TR8Ux7CaGX4C3WTASC
Mkc/G+GTQNmfqInlaSNMy2KfV2hIvapcptDThYn+FZiAzSMrzQQSdeBRkZ+ywDac
gS8eX92pUVuEuW2ZSfTpRjzX4cBmeYfV2aDRhPVvBz94/IA0bZsa+YRFVn+WaQZL
mbmQ4WjEMO0fKALvosPBvcilY7SoFCYNuuwe33vC0vUdobaWiUw+fvvg+jLkeZeX
ivxbNlV6OqOtTwzx+lSbe9zybT96NA1IsN0AXUWpAa9o8A9YT4zawlMatNkE1G+t
fOeDoo8bjtmq65hBHvA049Tne33UhrkqdQvdaVCFJNa1b7VHi7o7ikjilYbM38CX
0DSLAjwLUYJoBEO85kFcUjqVshbk2QNMCRJjrnKamrIdNsJnnPlxsIvT/v+IC5pw
acIB3RERnpg2Uh0IE9SHzecyIz757OBgYV7icdGGMli748Uwzd//S0JSjVsXbkwO
8L+JwpMv1dW0hxx9cNcEBNOr1Ek0bixAzJQNhocOBblwKTlMat34gaq4/7mIhbEN
xEZnt4vGhY+dumvv8VhQ+MxOCQQkiNrba1T9it/ZLR2/uo8BhhHa1jwP/0DvEwvI
seU5rMW46ZTIGAEIkYntL/JGtgsuOVln0dWy7My3nxBGbjcWBMoAWWgd1yVFJwRL
O15zzeG9D+2vgUkX/lHSrlN0Jpuxbl+23bZ4L1nsG/l13sVUa+sHTq7Jmy/Va/I0
8xMXfhE+QzSPQhowKAtwL2tg8qS06zvjUZm5c/Obo9aCfydq169DdHMRkWJgO+H5
8kAIT1BfmdwTRkmZ9IcEePIHxPVnxSFwzDI0NDLn0oGp76hITO7kUVqOJC40fpUi
faXaYNb7ZhVuDDAzwkK9lhiCU5PyquO+yjDnmkF2rB9uj3kxqdvvVy7sZCn4TH9b
PNB4kBPS/QnGPiAZ/AiSeV+PlAKHZ7tTpqmwojbd63thxOIqFWzOdWC6qA79e3yI
AppqEHK01I1ZFGGMYPg4A6fBPfvpBWvlOCIKF0ZmwYw69bmVVV510I5xJPq8XM4i
FH5nNtgZnBwfxJr73szJsHxfN9ssu8XTnhpFSmc/7KrZPd0I43mXriKBhPKqc+zL
/PJEpJh6B2pbU273W/wWILpU2/nLNjnbHj98ZUy9BW2Nep72yIPLWngJTywsQxB+
ycwWjMqu6DkDqPnpgVMmhDAKLd7cDzbYMnSgG7Ri64F7nOfbH1Rl3luBDeDzKav5
N2k43THQIMmn43vhdt5VY9SwKj/g2HVYorDa1OHmGR684zmo7sJQe6Bjrox9yQNA
yeuPquOZq0kZzj/N61H0udzVRLHqDC2RrhHPoJLzJhELLnroZzBg5WmhuGhzGzjh
0qFWaG4VRubQ80SDqq7kVR4Mxfjs5ks8Di8DaxakAPVvvrds/0Wtmy5OTXx1ChgY
v9/4mcTt7PrJphO+dAJrwcucsMRk7/Pj5dw8tyOyOWNL85ooKtoPuYGDqQxDuENF
2zmRpIzzAbqFT4m8bz/tHr7IN2IOtTjmt+YImyZFJQDB/6eCW+VDjcL1pNrzpNop
uOmJGJ62BbJuE3R3T5Du2GaEb/EWRQRVUzKUYTAOMyoAiFw2DGiEoSU/LBqF5vLl
/MqT1RdqWO7bXNK4Hxz45MMyNRzhb9aW/BWh1N66UmxMZYnySJxcvD4MbhscLKPQ
Z279JTbirhHsHxFYxg+birGOxPmG05vyKxUJFNhxxunDWCIBsLnn1yPI/IilbZbE
eb9lplnwZu2ZNR//qttUN5YZGrlPHV4MDFCNCF2imxksg6SpH0iyUaKbmuyK1Qze
NajGSqsfOxYrVPmMAQprni49GJToGCxXfCGssen3Z4ZOcJ8AJ9SIBlwkSsqv2IN9
5/BFAZuTb/eyGsWQxm8w58tBCEj5HhwRiFxhaJagxQmxETGaQ0Qy1J/vLqZvhDZ0
YPmEq8v9vbdLEYZ/VByxEjjCjrJ/C6zbAeFWp3IY6p/pcaStd/Xj98ZcLrwKNhFs
Hs6fB2xY0SB9OzMiGB5sc5PF7SDu+FmRnXnwqDyCYTa1bl1MrFh+rgNoq0BvUBZr
jgxjV8iaht58AjrsfvLCaQkZZq8PSK81YYtne9tQY3tY8i1qeE/8NBcrRKAAhvC/
0g+83UeHUzop0smajE+xcFq8T9CT3krFEnSQisIxUIoRiDS1HuA+ZRftPKBg4yI8
TcYr1gC498HQmeJdv6BWPjy46hjiG95Vr6SvB0GI2E6S4hu1BwMYP4jNCpZqLwsc
hqrhixJoXzfeNcCXmfHwcg14nRj696Gocbz0JErmp54OxETFYxFjOWloCp05nwBp
Nu8WL3p5gklPzvtAZosgC30WbVuMa/04OpfHOS2bt1DLk+wQT1SyE/ZpdxUG5i0L
Ju6UhZjTBCKqCCYGgKwKGgo3DBGIZ6jGAonCrMp7xYoy1NukRxGz16JUAcW49H7y
0qaQGJqAD6x7jUMiq4SUDs/VdzZ8p2KtxMqKPHOoZtf2DjZZlCvC8s2rm2lCOmY9
u/toFt4nsRxUdFw8L22DUQH1jEHfTNIpmfEdgp9cFBYq2NxCqrdlgGmlFFDn7nj2
DnDaE98/LIQZacKWEf8zCTUivSTBgy1QK/GSlh75/GzfBTr/YuPINnajhV7X5Y4c
c289PmEFnC9WV8hzpk0ytqPCwn8NMNwuUxNq/8r8znfY58ELpVzeSXjEeUqe0caL
r4+/fQgUILJ54Td9xnuuYHQvQ1FOWJfwx9yGxqGJqO3y5f4rm9ML3UexrI3uW8np
GGmuQ8V+53ld3AmiobtcMX4fzQHONXCMtSaC6bkcue9Oo7EZJq/gxmTmJGiQ0hyK
4qGpu3Tj3tKqRa/8XTFs2779LEiG8wmWG2NTVQIefbC0XdRjvIgLXoIm4rnQ34VV
ShT4pMiMlz7quh6Oed3yMm3q5WMRzYwDEn3TE0msLuda1HF9QHZ9gKyfoXRrR/rQ
C/l444Ob+JELKue2g1qiwZczrTm3FWuA47zAem/vhf9otAE/7lUfDt5VVf8+YDqH
A1QeMEhV0KdrRiji73zXMOt7QTBlgLu3ic7SKMcbLIGxgE4mBBXnBKJCjcVSW8kC
PkLx7x2My4KM5HK+Hu9FNUGPTaquLfl5wB/3AvAh1lAkNv2l9yktpm8TXo0jfnuJ
+JTpX5M33SU1JO8UlDe/jPPRJiN3Dd+rv82kzR12bDk99vzxw8TIM1CGHpTd3wwR
5e30CixD64JsHSD0VhzogenhR53Etn5eIN6T3ZuPvtvyJR3+mGfyNObXMJ9EC0Ki
GasXsr8Q3I+ClBv+Nb/+VHIxUtBZ4wnCHhsvEOD2p90Ht3yHey71T2XP3r0f0p3x
2gmK/isv6gtIZ8uk5fO4ZjxpVajaJ+buGpVz7FR2qH4l8eXwWZksfFtlcOeqIfHv
D+6vBBxsNouHeD4qneFALDQBAZ6JuYGHxelo+zfJpJRmkckmcPeBpej+8S2TC/gG
jURBiLAsY+CxGuBPDk9zBqxRocV88w+E+XMiszSUS5FkrUAJw9WuLhOwnwY9YNKd
OLXNoNVERe9u55MLDhhexvJDbYctonYh6MUFchG9rjVmp46ILoOBs6axzHCU+hje
JaJXo5IVFmiybrN6anIQtdMBlFDOMXWPWEEnshNsY9G/N4b5FVuS4szuyZ7+hxWD
KkmuI1Uwv3VDRZKs6CuJmWAIei9UaM4gP8azZD6S0jplhewy3HyExdr6rg/yX+Ax
qge5IQycE7ZLEeMA01ExXSHA8xfUKAqGsgOUY3XGOtBWOH12kRxcUfPjLS78H3qU
nE7EisQrNfzo1zRmk8/CIQglU5QyYs0dCYU4V728VtKrOv4sRp4pV29505GHTipc
CJNBygDuWa4q3vi2sWztMnagAQerRlnLcp9q9FJuuLHfWBq2qfopgVRa9oXjW1vr
M7UjhHIC387TWWj0S4A8zwlzcxI2AwthBABJI/fqmtamRxzWNGo25IukbytGJf06
Q8uVwrh9X2Vd6XoirWW9ZYWay1DxBmcobHl9Z5mj0K+IGg9pIVJM73p8sP9d5SzW
BM8s5Bz8dJG3eftb/weS8yC4tTIP8GdCKdgZDay7bR3Zu4vuCkNcd3QAyyO3QVCv
OXBt1Ayc6GXV8pt254s/EMafqXH/ZyTeA4odFdGVjcqyCy22hZdbyjCegUcIVQIf
ashMIhlmzzcVnRA9Pre4d2XfRlpITWQgEr4xaUp0dUs=
`protect END_PROTECTED
