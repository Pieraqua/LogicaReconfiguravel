`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ha5OYiTr5ICLBy+c5BxSxf63hxL5KWrwzzUO3gPkJNMiqBs15QDkb4XeraulUihd
rHS85iwAV4zKQIRsB/yTaDy4Twd95m+DmD9mkAiP0vqN+4fHwZ486RT8Tf6yMps2
fA0yaq3HnllKZZO6aYWLM0ezKgpEBD9++hBER6JmZwcsl/MgVUMuXD3onXoGc0Xm
Xc9bVXaz8K8clDDr3Y+Hm7ea2VD+oxFuD/lnzX157pfZJF30tjKqJOUXwDXI0qot
54PhDu03+m5Jhd5ONeZM4g8SP3AdVGgDT4TIa1pk5Epc0+49ZD71YT4ogLioNnvM
RTy5xB2T6qFE5VBvO4BYO8vvDK+J2J/d0qml9Xhbb03lYBbUivgRQCXYl5Xn+tpx
EKCEw1RscDfSYYTToE3OC3T/PNe7mazc/3j30A7NBRad/jG7OJxZtJ24gk/dhvHX
KsFwoLXzkG+wVNsMaDwH/fRftId8JdkJp+Ms1BbF7lT+0L8vI/Q53NulfDXnwaov
ZQ3WKQ0ga48Sd1i3BeNRPf2hxgxOQ7LlbvrKxH3X6b3Ea2mKWDMcRalMKldiDe9B
YHSinH00TDRURgAE8QflBPg9UrTHpZ30BzDPPmZbZxSIHj1rAA6bAKuQxWVSsbSO
0nfqXCGJVk86GuUmnGuauiYIG4WuflG3pH1iyPm3VuZ3jAQ0mCc+YlRfKq9jSvea
4WXnY9/9yEzoUcPnp2+aOC0it6bHCDvv/CqkZs8kZknReR8iKXwTM7Eko18RPj+j
L6F1uFaeLTT2aUdRIRdj1HI+PWYwqk5htdCslGNX/I+ZUeygOyvaLjU7Rz7aPITp
HcDIXlDLT6KbZP3lN2YiaKHx191nPfKDJ7CaYenU6gALpqwhGA4g55piW+Zt5J3x
6t4EzyMOOkL9bcl6bvXfMKv+na+dXT0D+6vB7EnCyjswL7VpOeztmmEWBm39tojy
8G5ItgXE9UAk2LMDT/pYNFqDXmxbwFC9MYMR2XjFb85Lmb8+S45zSWJEIDmrsFia
+BUs7+jchMjiOciw0+SyQ5NoCdUb1zpUqC6InIQm3WWGyAw6e1OQ3I+8d8FeW4fg
Tf8oSbzrC3i3gv9waDcgXWSp01Ldz2Q9brVHyC15gpH6uTp38+cUQrDzPmd5/pr3
Z714ZwNmYWytY1pG75Q7SVK1cq7ikht/hgWVAL5O1bS6N9XWhKsGkMj0O9zIeiUK
rriZEbZic8yGUan/G1VfWH2WtYoMahvhQ77nLlAsLPIuB+334O1eOqVlXqLvwyj4
zaRnMGckPBqpkEuC2YK7fd7i39C5nbyCb8OA8yzswzZ5uIyMK1XU6LC2eC9vgqqM
hKZE33QJCTze1x/2vsi5gsyYBRe3ERpdd5k9gDy9zLWwfazkeYoONzD7eujx25xh
NgH3OyQ5MHX3wjYOd7PZnDJhzNSqDu2CwxNPcd98VmgoJqBnQkV9kDTHTBBesc0r
i29g/QZrAi+R2VmAuun5mKhXnTcXHSgie1bnvPO6NcGQ5AVxvcNnA8b90x2T2H11
XYmW4MBwCMUIkQ8piu06e5heW9pGvg9JtWmK1JTcFfBxpLnJ0Bet+dw2CRwEMsIw
eOTzEhCQTlEANn+Je1iZVxYsatAQNR4LP800zf1+Q63gBKOuUjO/M5te4isJmqOO
usLqMQKzTx+YDG43Gxx0G5mEyQS1XbLfOj7Qll1mQo33Zo1fOoZ4bnexT/woXPDY
o1Eumqi7Wxqv6HtlJVDWKczE45LxxUNdp3U0XwGUP/yBB1nyynKiVRpsq0jdojLi
9lVmQ/pQvjNzzjJJti3QMqorN1ORRUaUICQDCsdPZ+4ERS0BqtpxppYyRzC322zB
HowqUyAmVcYkHn0kO7xXJXqvGcEF6ZYLWvqQ6j/wq4YDIgF9IEk1IqMEPUhRG1vb
CZyJGOQJi3IWq/HIjmU4Tsausqv6eUXAHVlczyViuMvdmu1KFOUR5C8lRhc5sXny
2+ejxuJT6BlUkHQReoI67Wyue+nEtIqCcB+WTevYYJk5zIYK8QUVFUax+VjruQVa
4qxEE5Qto0L81bUf4fd0cYqaVSoHDZHoCdK/F0/rnPfCoJamMV9l7gkT4wSjxaYv
D3UkCsHXSqdhMzU77y3CFFWLnj3MT1NDieq6uHhjNu+jahzAaJ1t47LtWaeWoTLL
emihLahEkbonO82JQ+mLIJBxLCBb0+2M8dE0zixbRnOGqufw59ps5pZEtaQ1RZjF
qUAfMp/GmUTzhdhuGVdENw==
`protect END_PROTECTED
