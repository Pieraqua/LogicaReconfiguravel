`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1DcDIl0v45xsYgdmgR4FBNLJAqtXqFsE+Okf6u14Ey7kWXk4iposXwrW5VaoYBVx
XdZ6Cx6ao6fE+9i9KsvhMwYKPRRI9W731925fkc60hChu1COV8SC580WVHJBZ9pD
ALh/zQEc9iM3nrH6ljzaboRNl1Gyhk+gcy3rpRioN58d8XX3JzGl8FLwpAJIPJk7
/fPuuYgv1lpGrJ1kakaOywhQXINyzrOyZ2WRhcBhvNnr+tFuCOxeuNeRjk5yQdrt
zDqp3EkrOObCAKaC0leOJbNpRY4BmK5StcqeRYi8I9gBuzWckoBMOoaCvC/abVQO
mvxBqAy3u+iumOA+iynqBvDo1BLoMh9qjmMbAqdnoKbHkKEIO0JGWXIn7R8sQX1f
9HLMcmLrwKz3B+yJ+5NwzYsbEJA3Y9VlLXa1u/SV0zurwklCU/Rr+6UnW4dz5/fz
X+a6o1mHIZydl4jiwB4gW9pa6py+qXHjAGZbqW32m8Lif5tNGFJkDZDe9tNxL2dq
q61zPQDP+DERqQm535eKJJoUs/NjxYgVYvkxtoE6D045JwyetLcvId15NFBJuLJM
hZ5VZrYSiI60hmbFtNY0v270VyMIcPsmpnNEmJoy3ye1RXUtr9Q6pT3Aze2rAlG9
Y5SNAtudy8ccWeI3BddhPI76No6OBxpyhUbB91hZ3TkHUH0mTh++L/SRJQ0x405i
5/ejdVCBXJNzo670UdFSkR2A9XrLXRrISYMF5KdxbAU=
`protect END_PROTECTED
