`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zu6X1e2zErino0zSdxH2+9FPxiOzoL3aEQhY3xTtqihAsBbE36HY92WxuPhjZVi9
C2iEpVjNc9ef/edH4gkKhjElk5yIgQmAc2SoM8rBzm6WmyqVRG2jQKc87kkgvruX
6v00CMof7Bq6t/hFEiNHdAK8dJ/8edr9Wau0mJ/klFqQ1NetsjaB5mBkahdx6l6n
1w8AhTZsP3rZUJAoMAJLBYnr/IEvNtm920rOOS6qJQdU08jJtcEXkn3QiPgw5T95
LVw7zktrgD9dGi2mUZrHGG13Sde/WrX7IFiUGO09cw6nq0epoAR0dlcxLklhOKcX
MJvB88lG5gkE9W5aCdSOg6ghQLBnDFFBMnfoRaFAPziB3Y8UVtlx5oGqsQ/u/Xiy
ebyrrLC9AgGnodt3huyvqwWUMmJPgGUXkEbbe3yksZNVDQYA2FrGIn7r3xwLYL0l
w3+idhwljMhmsvNb0TX+Di5ick7EYGpUesTeG+V+X9HSBTe+n8dfp4KHGtac824j
jbFyo3d9bmpI7zbmPAytxfbW2dUpQJGhmd1PF72+TVJjYt7xEIDLrNpHUnMi4nsE
S6M9XRictmApu6GQto/qlG8o/C+xs7MMpXlK4zIY/wRHipTGCzftD+jql7NH6FUU
AWpVK5JGPRvzXswPO8CYc6WsbKOyiLnTZeaBNFgnw0WEX8n8HgWL1bBDD/1INOZs
3WPxgsBQsXElmryn9QBIqqjsfPovK1CZ2LvJaWlUjsJzkYyrDpW/P/i56EuwbElp
N+NWcsdt+SOr1v/xFibmJiQzoXyLpOP//EPmAc0nYmMYk9lUfNJCY5cvV9v6MSf0
iCnVUFNTOzjkeFNqHLkyoy411gMOhi6eoCPxRfgy2uPfaLi79CTLfNnWonBc4xaT
z5SBrCLSGzyxCgRuktgCLhwd/TohGVuL5SQLDN7qmi22vvgpkDFWCjyoF9jJjgel
aJwbEgxB7iq94I0uNoiUK/Hs4O8xdHYxLWEP0Y21nG9DNzCvgMlGjhRmicH3l5pG
xc1Vz4jFszxb51ui3TQXW1WZ7mNrPq3PwkS3Tu2sFkiwLacOkixOSr3qheybQ/Id
S3L3T+ABaiiFQcSeTzC16KKKaHiQE/nXVPsqtzcjiBd7U1QwsV1h8NbudJS/qm3V
lbrUkaqCbHjtjOEWmsCTPZ4jVarZprdGxaZslfzFeidlNG9ZVJWYPQv3CqtKyJ10
yGuumz54LT30VRpj8eUbYHMOPwJjFUrajkZ56F75LUbOdNhcP/IYDjorfVjgxXuE
okd6St9F3HdZR/RrRJLyG1zpPO1dutkrsIBupPZsiUHKLZAz+QCPKhEvzWvyWkJE
Rp+cnz1Sim3/7TgnLFU0Y6i8uVrJQkNK5tb7pskqy58BI5FC2XWQTawBBqbWHtgt
5ZDP/DhEQch+cdRdQdV4n4DiAblMZmryDbR/kPxTbWnFUy/AwzcyUdUPzX9k74S2
MhJ9oJtqfnenCTkE6r9b/8bPmzLeeFB/3Aj0j6QZxG71cYWH93Ynlp3gLpy7Jx5S
zZ4CALIue6WNK4lWcOTRTWOFfvgM/jRzSMiJGxUjRd/0B+d3pWee29WGq3aX97d3
z7e665u9vrXenJMNdHmZVAYbBEhssX7FDyU/sN6MtiyTFU/FdTBiJDjuZyqfjL6e
jHVLqJEWcpLdABuP8/CumydlPTNnNBAxakV2ghxjPU06iNcHdGU9p9sfm/X8NUHe
l41QGxGnGkgoma0pEX26/UKnnGHsW/oxsWqRQVg1Gl/DHt3iEplXO+WYQ+VyEel4
CzlCU2Utp/FLDuGbhG4YS6oK1SkhI1JlpN0hPthjCq3uASeUK5Kp802lToYq36P7
1soy7E/EAPRF7RFdd+1PeCtSIfs2rn5gaYf69LilAHrVBvMWi9Ghd2UBA2OEtk4x
i1nlOHMzSVJbNjttBM0kud4DprrLgjcDQqbY5ktk13QhbduuZ+Fw/385goGO/YXL
sZCD0p65M12GDpQ/Q4faOCXoKT/tzHu9uQT42XbYI38LctehTdId5v5L5Iwi/CW7
VJpJRjiD+lNXErckkGcXSxDLVYGjOq2eTJeGchKAfUdOXIEUay9nnk1EGG7D1XwE
bnm3+kxS9WYw/XeiXUIc53i5jUMy3cQnXDkrPQ31POLTgM9ZY6FnWtWUIOW7QkAz
aZvjH0MJith9dAfhx3Eos9D17lHmwRJ3p/MO/AFHbohrptLoPRqPCKG5TMlOGG2s
9d5HnmvKZyF20dZhwT1SfKgP0SLAwdAigoK9pZOmkj2GcwZUFIS+1Ms9DpczF5Vn
BalTVGwLVmbwKfQcN/h3ns5wSbLc7wMqMt943WRN7dKvqS5yBe7d8lRnjXqZ9mmh
qERQIu9dmnLQ9SsfjjEIMm5i5PGgjmZxPj5ZBaVCuLiTgsnbrL2lhtaXMVMr/yiR
kBv5PhdAtImF44Cqb1CSALd9vssllmfSYUUXE7HStJnxEnP7QR7HIdPy2URIYS6i
YF3KmibLt/Ozl3Xv9puccTR+qaCYSqA4XatcJeNhA9X4z9wLMaupm8h+W+E1wlLn
c1HczfADWwlrl/qQeDlL43Q9ECS2E1CRUDui5jO2mNV0260BWDl0Nr9h+LnTXQL0
+8MSQXnTZiRo+YLPxbKz8X+ZVLdWukMfEpfqk7mOIWxDyc3ZdLHfyvtK5BoVS0Vy
FTS80PfVViWXd12klBM1QuFqOaVe5s89GRBEA4UxGoKlXiXOvTayKSv+NpxQg02P
oqH+qbt+6qCcGxbj3OtzYnY7JkTIsYND1frkXvzTKMmBiBMRDPPJcfTHUAkmaQWw
epfAbnokSwyXaVGlrH2bOzDs1su2+EIAxJg4k7aYsz22JoDHepSqd5Ak5MkLccAa
pLBvRAy8zQ/9V12OtwkVXArcYOMuAR6xyOoE1jMQxyRWhyFgF4ujPyiv8EhXEeQF
slcSSCU3wZFAhTE8Erc+JmQQrTLWLDVBbo+WdhtClow9aH9mbFF7tiOkIS8C1WYF
aUHeVHUdZ1Hny6pjSdrKOvPyk3/xlwpX2giYL14mKDbBiKTrZfSx04xt+q2PabJc
qO8/2X/bFACB22aubd/+mqVy6EP5dqhizc7k5ZbPaY8qmEiseakcgCcrXfz6kCIx
j1dY3rFkU9ms4x/WHL9VX9Ld5IFnmu7fB/+JVgtOCsaGx9ASOcltXIetNXzB+bI9
cznZNEWw4xUFW2HMK5JgmVPpp8JsE8AJk7KoFx4l7RzVTw4QxNMvrQpuhQe51hl6
OS0UACsRXXBs8k5TIwgPX1GAm+6A6IWgY50C3X6g4+7dBQa4E6WgHe3ugBsj0IrP
2kTnWQd93Yzmj/L8R8OsJdovmiNRc4O3HHOl7JY6u9Uk+jEgMDPDWj+MLe6Z4Cc7
qZICxFeOrerT93mDSzF4yXoHhw0AmD3tIvJcX15HP+XQ4Zux9aCm/Y9A1B3j3NQ5
0+CfOQ282Xrh9WqYrVwzC04UkRE0fTXAJTDsvbvJ4zg+eiGT5xAMTmDSQuiBxwW2
RtWWu5WMPAKdpJSnN7xGTais+JMgOCOnhbm2xD4vhFZaMw2to2bxIjYmYQSL4xkn
YjaBgKlB4b8Gs4pijHIR3lIyWA7XlJ17Per0xcRMEGpZb6xUFVose6u/QHsIADgZ
NZUD7jeeooP2TBDHpIZW/6OvLs48F/4+vykdKXNp6SQJhi4AmJLlFLeHJEqKlSDc
ppEC5y8Nqc5mlYCbdi0mg/vpKZpK/izlhOIQDG3ROI8Ga1wFuNIV4NmdxQCoEP4r
imWW84N1Qpn8++B2lo+Mt3rYIdPRdIl0LfEWeAQjZs2eEOUJktldMQ0ANUwGy9dz
G9QHc3mxpPVYeAGxIWew/TSJulE3mvC+TRDPvxqAUQ/IIRG+wIZfxp50jj8OcceT
MhiLAXg8Pip1rSEJE1SBGR4xLlKo4Um3uwWRjImSyFGIj5TNpm4tOJKOuBJ+xJ90
fKsl+7VyrL3wdMpbTjZsXNKudWtB7C+HfAOxg9T7+5tb14TQtj3R0rcu7qmdSkH0
5Ypza/se1PcYMydRc33u4qSenMJ/N3zWRF55+hU/ldr9rfQdLcGuhm5uENySU8s5
YlNrvTEJclWmZrbvg5TzkExXRAkvWgMiFuEf7c8WznV/TiM+Z6pA8l+1AJ5CBj3v
MR6YnofigEVlOzQ2jNSLZxOC1Zg7REa43alP2+bALREsk7YFnWu9HzzY9XhMyrWo
JtaZqjVw1TPYW7SLrOcjbLNybRHIvtoC0WDdN8k2lAQ4ypaAxYFIyQ2fVFh/OX1M
3o+L56JTrKj5d/b3Sw5eEjypCBiGD2q+3QK2O21qEBDldDV4I52KRk+9fa7FWiXU
Nq8kmJj3k5pgLX1KOwYdVcbSD97mJTmwO+Q03req45PalEi6dVCKb6rRdDBIWrfY
s9Pb2smiQlWOor/HW5VoS5rfUhNsxMFHFRAGoZWYh4XcUOINo1eNaDH9R/ltofiK
IytXBoxY3VQekBgES5Z+KrGR0x4ju9T4OJztfoj2ZHMN2WzDKpLjmoOCLELHYl1F
DUi0jcyXHkmXtKBHhlk96Bo3Fp67mmgWbve98xaxJYzzkLbbJKjoIEjKzLx8jHX4
cLV6DjLEd6zFJKsKn9kWEbDEoqSYMbuKISTf1pYEsKTa8kDRlZWz1w3AYQiWh6qy
52vrJdE4BBIOJFIGixiN4s7EE+uOhgQn+YPkP9F5q/hPVQwDL4V1BBnVTKC5kuXU
d/7Pd1lP8kqlkzN35kGSyLNwncC+Ajrcnjfd6et47JfWZ8Uz7iBYG82cdAqHP5Xs
cdqG2CfsJ2HMQqatAd0w2rHeF/cTbHkwFdkOBh1mj6C5RT4geZqjyuqI8rIh1OG3
geCayS7AL/IopuwB5WjC08UpMS2XsXdRnOaovDzoiy6vuQGTP8Wpgj0KAwY1covX
2TeAcqoM2oG/Gp2c8Lt6bAQDLw/oPWgS/Ewbd8EM8hoscVFsoj0ixkUAD7es8nuc
jYiV8t2ctwT4BeqpCBqZi543EBTvyRslY4/CjY4KdKj7m8j37k2i6mE5q/tCQXQy
r0VgiQhdxTDZYpzXibAn3o19OBk/BFDQleCt3E2s4qS/z5QFQyn7M6icYq99k1jW
JgFIgBckftA3bZ9UTikV1B0hvpFHyWZNmquTuLLvF40mg4qs3jwXC9Vb5FIESE+u
kQw4OzRLb1mYLNBNJdWjdzhmC5urcOmWqQBvIcRQ56EfVxN8Cm59sBMW6aN9B+5E
PERgYdAuTPuh16ntSDkyA+ocDQEEMMNNzhmqbJvoL/cqNCd4DuAJh6sI7v8px3KF
sV9kmn7N8IXFxaGYw038VBz6SVBlgDC8zJGuYPW/P23mnplUfDgJAOKhKWuu4v71
4rLelFfiuh6SMnqAsBhfIBoKRFrarZhwPq3Hss6dPy+W5pV6nrCrIC4yG5aoVig4
KYKP7Gn73OmK/ZKOTHhrS+z2V0yNLbqVviomh2CFQbAklWD4sdp3ij5xLth7TNe7
y5zagdyXxCSTvCWL+Pu0YZi941U1ppzIY8TUGShMtHhk3ftSf+qkbbIUxk+456X5
kAPabvNuCrdestrRymgVoC5dR2Llk7h4rNFZgvHlIdF/TntALIVvdkaM4cdjlObc
rwWgvxjCBVZdABWwVTjarxSbpei9B+FqS0UHD9HkfeNumO5BRXsi6Xo+kXZgTgMz
2P6pDUpYskItdrJVMppw+7GxPq40RkhkDZNPWpuCadocwupUv46jcAtjaPOgL15z
5H57oIZpKhoQ3+ZJNMehk5ZiTdy39Xhhlj3gSbmD1/lAponcpoJrCXeIO5wymzk5
Wt0lWl/iVaSb+nOmBl15PbscNNcfiK27WV/GsRg4Sg9/YZRy9iYbiMupSGDXkIKn
OM4b/yMvHvV9Cdu4lgfINm8JBrHoT9sdtCZeGMp6B0xaJOnsw6VkSJSsnDZ/Q5cQ
FEcgNA4PL0EkrdruV+hwXNPOD0fndy/FdS7RAeYJVN3jLGCtYdXtj0hv8RcClHNF
ZLbW9M+DtJDqk+59TCtt5+QYblXobGkM0oxrzkQFLYY=
`protect END_PROTECTED
