`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
glh4jooX4sQnNKLOUoRe+N2UYUMh7P6gT5jrAY8iQNjC1/zpJ7cmscx61swvh/T3
STdcgt8sK8Nhqp1UIX1PeLzycChF0UpK/qNc/T5U5nC/4caOmmaVCNwimM/R6mIw
Ff39aOUw31Qggz0EdDBezDwtQHy5bUS7zctVQKuJvBD/RNnvSaDTRNLK2NQcCHjW
JWmH+sEq2g7gRRLztLgMJBGIRQYqLXPK/tSCfDaqsKXUiVB/hT5wytGquSGKoeJS
NpDzVxYNe1KBQJvfuR+fvLmWqyI03/ayYZINr57xbZZej4FUhdFBrXHqHzjVvc62
0eF5XMHySLSKmn9ljLhPU3s5an3tAyJorTgbeUUCfj2poiS4IVN/4SRkXSSbinwa
WiQyX2fIKwidtFRgOypGBJqWLr2Ladzd/zIOqZfMGJl1O20YZNDLV6T9Q++4nKaN
bDRkpgdcn/UvvVyd3V/njQ8XIQibaVu4XRE+DtepqIYSq7C8ExUZbO1TBaEjufCO
PWhCsPdi99T2lNHv3hG2cLv3Xm7kwYhB+NHA05bnup/rDTgdWU4yPZmpRA9TBA6X
cEWO/nRasjKN12h+35dh308T4emrmxrdafFjbg15yzhVXSWTvVwkD5Er5ujRYxNF
zTMuxQvcSiGRbuSInWOCPBUhIOjjZyrADAh8S/VASGIl8Ppe0p1n9k9ZXvYnO5nD
beSLe0noEmhSv7djq3WVu7DfSB/SO/elZPrBIKlLszP+Z2N+sd18fjkuLH68XABl
nBz+VMl385BN1Faoc32+AHyVIs+vAMwzhWI5kb6zK6pqsAxIuE8f30YXlDE5bTIH
p2ijJmruJ4TnLPBc2otbnf2fILUxHOvm09Cpm/JSX/zf9KLCMOkh5B64PgDX2ObA
z97zY+4lxVOXgCTfJVyaNL3VIwkUsQT2YyNLQfqb0n3ACTEQASQtLRrtGCXbhGhr
SGJuadRmTVpYldA/5pmYhNYyDld8tVQZkphhl+u+l2oqcxCqqq8xEIV/viKUxbeS
7FlC7SAIDWgXd1mNY9bBzUD0tf9nTyeV3U1Y6kTQinZ+8t4tKpdD8A2lwZWVWl3H
d+CFUv9PvuJaOw57uHhjMFiCx/2belsl21IPZZQr8YpGynAbwJl9XPZcShdypqbK
2YdsyXjaC3vKyXvBAAO4zEPqrPut+BZ5dUJHxNA1LoMDPSxk843y0TQXvws5vlqq
7ONQqr6MuAi82pGXg3gHGKOM3GII4D8ofnk+DI2O1j7I3tTMCUDFWsmQUbzZuro0
CrzOqMOCwHtKG6k+/omaYGDMgJEnvzf37lbk0xGxnZCaELug9jWIpKFp/4c9zjNN
t4Hm0B9JlJHbKS3gQY6psREPnfygtwmQer5Z0tVvaxfmJecaVLizCVEk5mrZUSgi
WX/as7l+n7tn0oEXq7rHPSiJ5AUBD140oiZNEFauiJfqdVhZ7w92rjjEEpYf90CG
j5ibTxz4vTpaJt2KMYX3T7/Z3tt1PF57dPfJsHgkR9Cwm5tvgTjy0XVOPW6C7ocM
CcRbjMIu63adIreMQ4AlkOKN1uoAMGlk18fN75/bRmcrg/WMk51j1lxB6ehbYQV3
vehOF/zbtCgAljp57H905eYAaWWFOYrLYI2tHCjwkCPCWgrVriy11w5CiLlWskWD
vbMbXsaB8li0NRBKm39NPeLj0MeBJyVp5Ht9bnPPyn4oxyv+0e3YkXrQsPI7q3D9
/EUZYDD4a8DlMUgjzUGNZhzyNORCmhAJs7nuke+0PKIGbClRjiHIuAYxnm/Vcctj
`protect END_PROTECTED
