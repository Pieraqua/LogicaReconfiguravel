//__ACDS_USER_COMMENT__ (C) 2001-2022 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
//__ACDS_USER_COMMENT__ ACDS 21.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ltLyxeI5I1RJQ6AFf9WiA6c8E6kDHQszJ7CcvhcuiyYYcoeeDcHx5OcdsT5M20+bcn3VsJxrFCbr
JfynXsD49O35DpUZd7xiV8vIFf55KUGam6TXbwt/3CLlpmFrX/YXOPodTEbx17UKfTkW98KI/Ja/
ue5cgvGROJCAXzsA9xZda9NOpvECUtWRM2LPlUi3jMIedpE5DMX8fyDmkVqmdhti7eknza+/YJ+4
tZOJuIqw5/BJTf+3TFAK5a5BjDxPa6eSyI6IQ1lWevJYV2e7f2F7XOAk4AX4RMdwKR4JjlpkBEu0
rjH4oVD9aaaRmtQJsIQ8CWAPbRVvl16V3hVb5A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 12704)
O8a7YFFnRgJPK4B64n9z/CcoOG7iko1fImywLSLb3HVQXeJhTYExtLBULKHSoKXbaG0eInmxG2DE
pJtEjVEiTCYKhxTQxZDFAiY/aR9Zb13vnvHsGlsQXm9LVhVtOTjzfkAQiaM+6z4dz3oUCY2tYY/G
wcm0Azyj4EAZWTAf5570xWGpgsk5Ddfnw3uqaSy1zNgkRwZpb7r2IpT2hJCdXdliOKWGEMJyFj1o
mwZW05V3esi+pT5WpRuTYT7L0vJJYWkUbxniiWm5Rb3qYBTzQ9r1caV526SXJ3fNraebUiHyFWJz
tcfjK1qsAc1z64dGEGbDgAPmMBrAfiKahvBJFyYu4N+QQzHBnBDv29MCC1Zgr5jbbnSob2mABt+C
11JRGMUQCQUFoRnK5MbXrxbGkVth6/Bd88Ed5pcufMsTytlXRcMue1iZaJZXLoAfr9Tjal4+Xo0v
008BLIz/ORohuPm4C94OTwZqQPyquJ+YhtBOUFG7sF3zTnnsaJIhsEacidZiGWTj12ImwWTgPuLq
8YQMIKeWNYFZamBBilp9HhX5XqZwXo7brrT8KAdg55UvPcdLfwRLIUKdoAQcTrGhJ0FTL1UxPeit
wwLvsoa9ZZA8hLWgC6DylOVJw52sxs3iVDMjF0y7hZLMlRIv4TUgjkStxncVEyicHOJYWpaTubwv
qUG1eU3BhXUENCToh2dI3slQS68CYxAYg4ffOriksK4S/4e7G82FE34y769BDDZA16I2tShkWgcl
1UWIMcLvetWBsDFClGbWQo6RxmKRgKL3fnzUE8n+tcQxyt61XYA8QOzJxJkDvP+AUbh7YZDio3m7
Z2Uy0gcPon9ylhAQMvl1cFfePIbb4vrK+RA6wE2xcSDu9O5Z/c9B761e5gACWrDXg6150qqqioXt
V6toyhGoK7U+uwxUIPSR1XvMBB3cYHwTxDWioPJ50PyFMm9jGRJK6m7DCMBOM1iWjzG9c72OYAuU
PD+NcP/iSLtYGgCjG4bqfIu3pmngbjQsvEYlg4GZqiZnxdtEqmPhwaPO5QnGqyeAM5p+diFMx1fa
xqubs5tqztGlg2Rc8WreTWi1CxVez03st+EdrMOtm6jJtEh3LklQhLTaem5iJi+e3FxVMFxLkPDC
J2wesxhfH2WDLhy0VdWM0sNCWI6/wcadOcLjO/U869QFQkGEiBawv6Xq1dnFDry2BvTCarXakiz+
jJbRrArcNuMAU08qIbthdGa3ax3wR73TVjOjSx+rf4mB+k6hGlrlUGzSAaGtE80di3jYrC35BvYp
6SDK4K5MqqSklIuXVgwT+FT1utZJLL30GcxWY+r8Lq8dcsErPyr20VDBPBslKiXa19Gz2BxDlCmE
2MAMXp2+WHSYWIuA7pbGx/Y2eJ7XkLUVvNGWPZsSWSZYUL1s0sxeopc2jWXZJby7qcc6mEY04z+i
G5lzHVpsXHsIOwfz0bCr0ucCQYPqwHkZUCKxVqqm4juXQ+gc3sWYi8C2VegMUsKROqjEaHfD0oEu
p+OJG4XYJO4ZRT04nvE3uv87ufebWNG6gg/POCArgQ/MIL3LIJnf48BVqkCFfwPCueP8ndeJKbN3
7Fd+Z26/VwiunPuRHMtL+U4gFfoQ352fmlndPzLThCDUnHrZcQ4fEXhi/fqJvZZuMvIZcheEJU3C
VcNwZ1k7/VgmBnPvjfy71Yx4Pm0J/BlJkV7+jdNh0xMgVv6EvGE5HvMX+ZPeUpZdBqHrS69C6w45
Jl1lxw4Rls+Je7MQSTtGjvEZ3no6oVm2DOHPgCwGPCIftJxu0OYsm6DI3dHPcD/sEMnrPRJH1tCu
fKryfNm1A1MffSRT2ORYSlmX94/FcSowvpl0oT3phtscGi8xIZD6G5wDBtwT8n+KRvgozX+O+6+0
Vd/OANxKv+kDA0EMgi3FhiiTVYrMIB/lmqFH0eui7rxs+Q001/Vrh2X4SFMxjTYop9Y030/lnTIQ
CIGEMv0YqKOG/ya6LodMHtL9UUgSuEcbtAYDCZxo71o0+WCaqkhBPme/LbbWPdcmBrH7wUOxIgF6
tUwhW7XqKNLDRXEGIpol1H5nBt3flgwcKHRvxVOCCAGFW7QFtEdec6Q2GzpHTS+EhXNefNxwJkOj
ifR3WOOYrBPWeGkoCPbLIBKRlsBsEQSjTgUftlmzxVIhz8xewfbXNFn02SbmevrYB1TxyeA0Sv+f
rFQYwt2lsGOqQn8IfCtuVcFx54e9roD87CcifJzBw2WQUwl5aJDlmioY3vcLGmivMgeqxHkM9H4q
4NIEmxlPG42ISh7mSr/Cp73EGolu4m5xp2XwDyj7uv1YBfk5Olmidjr+bRaTH0BOOopHbJgv+rGj
KoByR185fHWen9TMd5NHgMs/SBIyn9E8EQVOoNl2Ubu07CKSWZoVD/jJh1D2c2hku7KHhYYJ1sEy
BeNkEQEExcgYGzTN8H9Bfg9JcBj56rnHXtQwLZETMmk+x5eUCQL7bbkJD0dEKxwiVT/zsCtZXzNU
qmNweKmIbnLK6QnGUi+Vn2UY3lnMAsStoJdn6gJnY0gOjHmvpDk+hbfVrk99Ro1UZrtWVrNuWxmY
0CS0GWp6ptq1dtHX6GfhIyaeKAORgK70ZH9xh8ViWWU8OVcRwep3BNc09AiPpl9SFRhIE3tWDvzo
Sj93+aE+J0bjzdGrmwJujrBOI5y2QuX7EXUcV1ifqa+xjwh+m0/TQRiBvwjsPEeSF9SjZY4zSSPv
1vmNL9mty5XX2d4aq3M4H11HVHoGdPIf+c2APyJZQHUfNzHGqQNWBuxSp4ZMi0L7/GhXq676bHYj
Qut77T9HCtBuj+/I/wapcp9Icuu+kT1XG4MkyOvXWy2HnsJ4mSEr1cDpkpmmvNym64OYHh/VmFx9
qThVg1paJTXcTlX3/hBRJ1TasrOyDSAwIlyUyPrGa9ndZW40HmG/CXBc6A46qdmCsghMDK/FRtQ6
CHZkondNsDwrKbSeBQ3qHtwhYKQSNWqVDphkb00g3GN5GNvF+imL7JWpvLz8NN5FLF2Ird6P34DR
JivDLxTpZPkbRlEK+85WKnTwcZG2tCLNl74lcHEAKTsQfESexT6leBklUZUPTxj0BEAILjHAQb1j
o8sxQA9fRxorGri8YdJeU+UmRe5dxiToA1aetVYTooWm2msatfcgmIb7uD/C1qXcxRzsvkdPfWr3
NVQPSJnDhuKd3hnQrbcX4bxrNBiy0ip+GqZShbsFqTKtIjKucATZoG/Xte4K/JiSjvJcVKk5ZyRJ
dMdszUHIOdETCgho52ks+LR8E/i+5p0ZKe1HOZ/UTCzV5FUTwZOSn6H56Lbyd202wKX2u9px3WYu
yB8HnodMuyNPnGdrIz15ykCqCgaBFrrIlJ/ycwvWCpcR5MN2+Ceyt8pX8sP1KU9BOS0NuK6N9Umd
MFFXDnm6N8qsabCA8MYfAF1+obApC1nIkjg7AVlJJPi3UNo3ugbBRevuuOO3Sv1ydaGftu4vyXZh
+Q6igSnNOHHhX5yIUsbyUddw7yxWUeTDHuajyccB3om6Ara0YdqltRJvZbx8lrJHcSSD7cdhIAMR
QcLYT9FWEs0M4ie1p8GxFeFGV9tzNYjOLq44DHpXwyQuq9Lg2AR5s5QmC/R2eaiuE0yJFst4KTaC
sDNFH5JifJE9a4uajzTkbTwKWEexvibsPIOgW7JaqVkntb/nY/2dv5XYP6lFGsB8myLlEF8lumAd
CbwIEU47PmbYIPqu9btcG/bhW7vIb/hsPwjHzaIiCvq4GxRHZEjo/l/ETc00zyvlhx3q0ruO7o+4
ta/vAlAE5h56+/JfX2NevCcCTRmEHzPKgETX7vi/BbYhTuv17r6dwCKW8BP99pO3bSUvzA0TOlzT
jqcT8s2ctS+aCiM+PL2LgakqY7l8YwbbUsoUtImYMYtIFcFkag75nZsPI/P46BoXaMqrkf7rvfl0
mpycH2ceAPepgfqNt5+U15WmLAquRFzAY1FpjMfQmn7ZN/K/J0dYiqBMJQRM56Bsith8evSprNj9
pSTocFzEMQ+FndWayt+cW8600BaIrVEMtb6dfWnoNcMzCAJRkYfyqR5fQWFAs/8yQeC43R02T3zb
mPd8uToBuGeoAIx3otq4ThojGmXLfTj99EKqwhUfIEz2sSE7Bk1B6XC11zDqJiLaRdpZqVt7+gtc
VXrh5EomuAPCpLS5rzxoOi0W2a3xIr+yzlFuepKrmAgB7TUOMZp09Oo+VsLaCJOsO5wluKuNm+ow
oAtOk0QB4w9k0zWbwfJdDHExwR6YKOzU0uWLVFJXjJA0AjU5XwNgA5uX/2NI+RrR/TuVuqIpU/LT
/CG7oug3JK8Gb82LdmZvbsMXvzSCRQb1F2jBmK6wd+zQY7kzKCYP7F0XyFISH8LuaA/vN72esQjW
Gz1PR1naOdUicKbPUE39FbOjYXpkF6TNI/mfg4yPdgypNmBkqhcrsmvjqJWmujnOuNIDceTnQUku
mZIL7oIK9KhMUIC/VhwsI+bOv5vf9dZM62VpAJ7qHE7B3gSyKJgFZtpOZyEAt0RsjtpncVViPa7b
wjxtDHzfFmALQ9KqVfgjFB15uAzV398Oh269UOLSUqJN8Pht3Nro0KDCsiieaKClx7J6CaWk3GUr
xxgEOqrEmbZto5jmFjQkaiLfG61xo/1z/1FPt52oqCPV7tptuNBj0jRdpvGPU1JM+3Cpuz2V0HQg
Ao3/8IgFZcAaxdB+n7FdsyrLckzoniVYvNa7XcGF/gvmkHYS2EOr6RVQDUToBdoxESm6X/6Lkzuy
XmgfjLe3kb9pIZ/0m/koLWXjcFYpJlZQ4CZFXhugg+Ot13yzdOa68NTNNxfbb70B8lyICxFPyokb
DiMhx3zfHoK+2xBCQpu9FZS+r+bklrHksV3wUx/x8NBbVidBHb4dd4iAgd9/TLkGbZQf0LgSiKhD
zfDarAZrXftc/H1IjUnt4DtoRqwfzffoV9q8QUzZICplu9jQd9WW0TY5bunqa81tSv7h+TnpZVJb
rgXuGrlc1KRfZ9Ss+COTQD7NoBDFIcslpdkUGkRCT/69FVJtqLmH8C9wt3ox1IxNXOCM2HgWO8NS
jorIi7htmE8jMCsBG7LEHM5Jmjl4Q/wYH1NjjaZKCA6p3bW1xW+S8+qPE9R6+sb5dutsQKhS0ZwO
q0HkaoNbfuW5bskcR6IBxd+BJBnSBEAHSrmEDms1e2spmszGzTgiorrdHJeFw4Nh3MfBztGwnSaT
HYVSDK2fN8OOZA2AnTDiuogB1nBK2JvPF6uto+eqH9QV2ee+tZEjmccV8aecV0NCQZ54VLnbdSaK
SchkekxZM42bNSi4T7pEe9wP4kyTLt1T9BSmFHj+cLrhzBoDECDTp6B5OfXGtDKBpXgOFfxESb9D
Alb1Fxyp4VxepNplL1OHEkHoT5oGMMBeTjzCQKWQrmp8VvruXptQkJlAvSBN/cE7wF1zv7VIvYSD
yYMOAR6iIyyBBfg1dzr14IZZZfCDyRlZ+h+Ix09ESdOfxX4pTsI1XhlC0fUA1dX/OWLjOw7egi3b
5omZ8nhOUj22VHrUqFJNeq6jHU8iKFJWbBQuNULqz0/v9HwCALpR4FmqOEqhcgzwEUQapUyBzHqR
XVWtsdo8IV+blMWMFsjbMjWAhgl7y9jIsEP3XYMZwRQnlQEB7+sS2yZU7Auuwh7D0P/bvOXJ2OgH
H7luJUI2cZKWJgmFMeZHwysCxkAXcz9DMF7MUX6EY4HSc4obY27pWbpHfc6lawvC1sJ8LWONeKI7
CjM7i1Oq4VIQZvKzO/tfmRYDBI82rDgM8egDVxAlLQXRzF6NFzBIYipaFowvWPJjAG85aEvVoxU5
e018adDvLmaY7v9sdJ2rI3vuOTHAqu88T1jklAFmcAdE0gjbeYpSV2S2yCCxYB4aNHTNgMu2OJ4R
gKHaWap4Y1MBs81UVJAU3l17E0BR57+m3WybtuoVd66i0rcJ9jz/rjHYIaChMW4xdoqDnKyFV3sz
I0Mwf0ERzgsaj0/6IWE4L8dDPcyDaxxJvhoE5likPUBDcspXFzGrukXhHNw/Mn0dB9walpgUmver
tpSpbZVr5Rm6iQU/hAMRSV/NbgI3vEmxQQ44gmKuSoVvGWRQU+eNOh83MkbC+hUfynSIDutNbqiu
XpqgD0BHuWzs9KYM/WiS8NnD9rz+Nxj98Ac8YfG2A2gSObsbdBDa2B929Vt3O7fBhJupMkuoK/Ly
38t6Lcy1ngEvOg9Nk9RjkfzvCdvCq0QiwA9d0UkY1dWJHx+d+t632baDe4LOxWta0BguYUM5+lg9
usky4QkbdcmpU2JoLYgEf6i2UZkJWy+s9qByzM5mG/SiB1I6rHQyjz3qCR/NWnvAEk8Hm/GWIqpg
cPivd0Mc9q0kX18TSp70NWVzlLYpFLhIXaJ2/XInelqG4ntKLJi6VVZT+aGayo6o8Re84ojcPBpt
9GKXSOiPjtoI35nptj9uGcFNeE84AjVSnkwko8Y9TqjzKfmLiT787yiUlfF1aWraadv+EthOEYVl
TcicTGIuYXB2f/RxcoOfZYgwMzUNEmKmb9lNAlyOaBAqHpuOunvqcGYiwto92MrPAXUIg22gMiB/
noixSKaTyqBAYDy4n7y3RZT7T3NE5cr+kunvNiUIwvUuaufg1KCbDSioKxEXw/ZUr5TptKSXKA07
xciqG68IiQbiRfK8qof1qLujpmwqDQtLohPu8xhixUghrU5oerFx62rMW4nKvZHgU/HBUzvd4Utu
th6Z16BN61pmR6YBIUOXdoCHGX2eO0Je8aFEWBw88cn2aIsAqzRN2C4FofhcKiRy4Vrt2hKYd1wk
N97N5LktKN3e3GTk3xe66OXRgjBDzmuZZbEc6l8pZAj79+QJRy6NQVqsTdPji1U0VvPhT3CjRnD+
SN/TwouxP4qllAIxEkzalcJZ2Y+zj04xivIcaZlOvYqF1IcEOwxOVmdSoKhyQqbf1RerPdGNjWRz
XV0MAyDHgzj5hcEssYY74IuhJO7kTMOFLh/FnGd9v6cvrEuB8+dxSvHH9bGqW12kIarV+0Y+zJpi
CC8AfpepT0Xt5TYfSmAqGj3sZ3Ua/0U+Gmn5CHiT/azDeTY2IuzkjHEsnWD5ozxkoRCjM0LyAQLb
Uzyn3DWBxc/FZsNL/tBH+3JOpL6QKWuR+/9D5b2tQHqCfpd2Okv4EPn9yWQPyBur433rZ/TvYz3s
maMzk9ET5u9mu2FyWb7IVLNbO47W1QWY3k9vnGQzLmZjodyiOUyz4KAe456SYZNisq9xRay4qjn3
lWl3Ar1IlBTw4kq00iEXAxHK9wnv3hxsYvjFdegY0HazKMDLte/jdX1Tz5nsyP1pnuTHwrboIJ7Z
EYIh3RcAGxv/lp29cJujgxzRHfC0Drzz6zC8TCN812GS7h8XQAF9UJk3RoXLEzRYjS1YiIR0BtPv
Tq3zjVUlVJvPK34FipiWjJRyIHTyVPVKvruGWxEL+hrlDnSUb5Y2fj/Grn5GPCbT8lCERdem/sVB
tgE17+wxj3izqhaFJB+VMNaAXkro4R2/R+pp1USJ8w3fwvsjt2rv6sYBVqgLu7rThouBrTJZ9+41
LFjjbGOywRdnds7iaTngsvKrqRsW1tnlN70DLVGnBYnHJtILUaXtTt5WaISA7gVqGbipr+xBxpox
lvWqMRDBaiv4z6/Eh3kxnUiEfgRg8mT3EWBGQ5wr+eg1r/GjqCvbwujDh52pFL9rpfCAP9B4zwhm
9SMzXIx8erPPj+NfQu2oMu3OxF1JaN+jXTraqvXKLZktICg3FYq5c5TcZv6/7nRXmaGCBp82TdAL
/FiG1JTWyL7sZf+MuE/cC+k3NA1P+4KkZ2tp+5LA8FvnrAhGvy9od9WNCXVugw2ekfiVnf/tidZC
VvalGgYC7MXLszgegYXmhaoGKOD3ew4sqzjEsh8aWoSVFAmz9Lehd12AquxEWJa3pwDNTrXWIStS
6iVnZ7OaDXcHvthUMmtkgsMH8x1Qmw7HRHebJZ24OznzTPoPe2cR0SBYUEZq7TVVXNUNBrPQ+Ghi
CfvP3yXutxGa5LkaTMCmR2H8NK66GezXfXvkrU6w/E4v3dwYp/x8plygI0ntr5RYPr56GggPRPqs
5nP7ES6Gxu1gYuurGcRe1RCVxHleWu/8juo7IvrlDhWm5cGgFLPXsPsYMY+5mcJOb7/8jAMG+d5X
3QSll3WcsZDtNJ2t/Xee9bRrksBvefGEKYWQBCfxKAs8XGPaXsWcQseZ9X3WH/TOwx0Ws9B1qxdG
fh5T9ToJEcdzuABwoWW4u7ev8MOmGLMWWcsXUjP7nL0IWz3Ky5Hd/W/VyntRG2eXiYyJn84+4uuI
kHuIxDMsA11TGHE27UpW1duLm3f5IAnnvTAdWns2bef4GSLk1+jChfid08oiUmivzdBosD29OKZo
XHjTNTm2Ba76OW1jA9jZKXBOLxBlm2AAnFJVYobUr+GSr/Jvju/MDO+P3kGvauVOZOPQDaQLWEPM
Cj77wY2XpX5yv4vAn3mKqqbuKo9gEV1MfvHJITJqj5jzX2MhF2HI6KbVsAGVdfmZ7IapqI8nq+9t
VLsbfCDtadzf0cZQQWoKAQpzLwZeFPW4ZJOwxQvw179V3pcv6+VDaaDPCTKgtShcJBPb4heecfvw
Ut37+kZOGuNKOyrGazNxOqN6AYTPz/ARjKVO0jgCnkR599OdbMHTyK/ouDnzoGlRnUnhi4SYBwjn
otfqcZpWuUD6myRjE8LXj3zI4z/ppXWpwMhRyrFRJiB9gqrYM8fLYQIo/+ynzPIomByM7bYFRgsI
ASlqXqv7zaa9U2u8YyMqfQv5o6/xJch1zBNpfUrDXdVTg7sfSoIaSLpqcEVRHmJZCpwGatpOcDyq
fXuJqBnN1I8X76PLiNNXgjyLUmsCNThUl0dvrpv+oyxwZ0hE9Tmo+PCfriRkrwJ58R6cGtXMGNlE
VWujXtI8QT/CINuZvUHmM853XcRfHRysYdIZu0hi2eAVsB/XXMndHDGZpSj9RLbpCh43Uv5Amh5U
TKBC5TNTg24/u1SmkuwvYzJA4uAVNpRSAWYXLxRBRoUOLva7toQut5ZsGeMEwGCcJFjUZyhJP8e0
uuSha9BE2bOgOuK0kK3KVKHWyI3oywUH4Syp8bAh4vF2WLqaiwklM52gXr/qFDKwW4c+yTPKqT9I
NVXlAaC/c4OnS95OiP01fbhIW9BWuzL0hdguoieCymT2ohvkWdFR3ReNFHRqJ4l+AUQLjrzXUjgk
ziggvAjODVeUxgeNWy7dHlOLURbo4sfpiiPo4Knz6LsvhQOoCkjgg5SaKmEJvrnJZHjHwzgcaA/c
Hu9XQfN5rdk0uVT2qR30Ni8hBKBsE4L51CA9VD7Ek4Lawvm0k6KFbuVbCPD1kv4znAWRhzZEWn9j
AOWCNEEj7bG+dyPT6g5rsTWxE8pALeHteyk2VIQO9p+9wLhJL7tLk6BKBJUD84H6IHEOu6HHkNwI
FFTgqyo3q6NaX2YeJXRvBY3kbGGtlhej4aNNwyOfLbBe1bA7bnDrJfpfRDN70nKpXG9xe1KrBJ+5
jRjGFzT7O4r4ccY4f/FUQTI4iCsQ5pIl/GotF5QaPHtX9mwoOPtMZsXhw+7V/ctwlbwBKafXU20d
cJvOuIwyQ/jAmRS4+KJTU7vaJH+5vcQnjX45gfLogQg+7HczmnNQ7O3Kz0XWwlQAISuWCzg1daGc
TJxcregXmwiiXN/wnRCaDuyugsQ6p18KeVNSekq0PcO/XW2gFzyv62zUjHEp8DFe9N7vUj02Cewz
Oye/Cg/Bfg6wWGaf8vCuUwCkrhjTtL10xvXn8MfflJL16IQkAue70eZDU0gvtQoZ8C6Ka3nEAjl6
ol7tLADln7mZc6a9o5FLbHWWoLqDHlGd++F5953KKa3t6etz3tpP4KfcnnMyXv1egpLnqMpGcCLZ
87ZviBEBTkU/9pQH47XBwh/FRynSoah6B10cEMPYnSbckgcZGQpCyUm3JKyjDVf9cxtSbeMf0hKK
b4wZyXoXr2v7w5meY8s6fbSOJ+v3nyISggq0nsw/E3uuQ/0kKQOVv+lIIgxtN7VKjNqxbVByTxlL
5yxbqMO2CsnQzqoZv0ZiQIuySJhpeWdxAfdd0a1JYdesYO651exwAgRmyyZBeRrA8sCwwo9WHLBu
0ZvyKqXpnQaPgpezZIXNGKh/CRg/mvEq/W2CuKGgttBIi9ZC5iChPUQfuECuIuuodDiY4SmrtITz
5eMbcnc1VdSHU4pAyZeczymz+UUKiqD9AfvuYro4ybZCY2co3QVZL/+EAM/N0o4AleSFgV83i/eb
2SdfGs5tOyixXmRevKWCOngMJXzdeYk6lHQ3dwcl4dJpmt/R3iiM8zpzWHJ6asWnAoI6JZ04r4+P
5pt1FrnIOLDogjeLFGz1TO8u6NEFtRplEUeBWnwyM+T/FZka3Y59FsX5HHBIIOpAVVjVeS3VA8rO
gd6PebAeaPyqKwMKCs0RN8arw3pzMMH9gBw/Ekp4T9+63VvrQ/AsAYeDpwv2hkX/btIh9P95RPlK
zxUVUjanuVr2H8hRTNpgHOtXVKFt+hHC3Tod7htMvaPUWfoE9yL2ubiHIykgLZytx7eqiqqvBJ/e
+VYy/AyDVEA+Wzbiu4rWNpOLBcUtne5pgLSOdtn5wwKQHrwCkue2l6MsNL/Anv11LWhPewixGxfh
b7AFwYZIh6ZdKYp+9Fwvp+MykBYsR3F0j6Tm7I+gKOzG1nQpvfng0KfZEt3Icr1b113ok9U+tRrF
Pb7Sv8uTFSHEgslX6kU8IYnbe4S+fiQKiSJjbrWiRKao1+dEN73qDzGRE+RG3QiZx6DlWLawHTWF
Vkk+8uyTsDwuqk10wvnGU+0fXnpm0iz2rpGaQskOd2ygvX6FOF6ifktI6MpfeK1FQuQAbdv4NZLE
IuGHcMxVcZoRgIT+TkuPOnLFIBW+QUhOBZVVmQB0A9jzcRD6ArYuxwrLXVWRe6RmPJqf22lrWXBi
19Dms953UQKs7P/k34MfzPLGb0XB17p41wSQiaJ7g/FS6CB0dhyD3mToZNZ/ajRMId6G1FTzaBXW
Q9USOVqxqENmTb7fgwck+tC5Ck2AVJZjWcZE/cFxo7dWejKDDb7ZRXUwUxYcZDQigQ4ON1wYU2I9
YTwzdm7MqsE0Zi008aDI7WM5IYLMB2NGr0Pmh3N8Y6olZKYX48HG396Hi3AYwMUfWy7a8Sntn8/4
vPVI4wJZewp1yNlwBUKNYD+fcdTorErad7E06/fUbTAzURw+PK6WEYw+BuoP7xXAQYCvl8+jLDT3
ZczLPraamFcvLinTAU2nT11V3DP/xZlPx8CNJcucgQyXrqeDifyWDUfQJzpuhyTgrCEPDtCYlMj4
8UaXglb6LgCjYggPPdiw2SdQm6asWiSP1pVnh1FvQ1B22Z+N+x7Kj6SXcnV2Lz5R+V4OVRvY2Cme
CJ6wbYDZVsjID6Kcx8KfQQb7Yuhsq7JEKQUgeg2p9xZau4l7tZadza3IV3hrXcN95AL62AtnEeI/
IjXB+xAHOwMAPmCI9OxNcgDGNMngvAK7KxFbyxgn91hnUhnvwyL/fVo0HL5aPQeVFGnCx55TLFco
irBSQRGDhxcfZb0bHyf3e98gz0u+VSSw2dwcdG9RQYUhniIYuXJ4WeRXyLZfpYvpmcmJEnpSpbwQ
LBenSLO/n++EOhGYlZDHo5CP9mR4YqWRHWWyjwVYRoWxY5MkuGBEDJxb54gJOBQ3fmjzyjfZYW10
0KY25MfPyDJRCTFVa9M6XljMzRTS5BJ7ahEJ6e55ZtaaEOcyNn98FwCAK78A/HIGTJSzQUseOgoQ
jV6tX0yLRPxt1FWsJCgixCqEj4NEYHFfbkXi5F//SlN3ZZ2/MAC9a6P4GfmAuoPSuqQfT2n+9U1Q
hf3blhXNDidIQQNtycMLzaCItnszjWakGyiIU/DyVo/XNY2/oGfbGJQ3Huqq7gGtQRVDUhwkyl0q
t1CKtCBTFZucOdFBde07LhvCWVu0Z6AULWDPUkui1Td9BWMg3gTyuZXo4y4mx8iSpInGHZnojlVn
qhhwhCGDh1ymDFE9LHBNGlH2zd1HqMy1aGVU5Nu4LPbfOzBKue8v0JQ+RDklLPDWQPKDT7bHZMbm
tA0QbPFja7rhbnCsOFq1bLW8DJ43MTZ356yxHQPjwzGK+L+7bS2UiCho6UgqLwg8OwSsTZGOTe88
UibvqABIQkCpQcTANXqbAp+vQS+3RQsfl/z5EihFZCWTmJxZISPPU+2gMO6bTwt7pp9Tv0GdgVZG
r1S1EyMaX9uxc0bVYDjFM943STt0+M4sVlu8C8R7JF7ZojlLdWsq4ybjiTpE0xJMGUF+mJqU8Qb3
hxC/3bMq+wYoWgI6ctlJ1Yk08hyR6mt8mckhoLrwIED7MN3XwIMhYEt4L3o7LseQa7QrJ9LmKO0M
j8Li1MqXLm5uGYuDhqfS5lsmPT5swZsmwh9wR3uqryzzpExlmtsyKjlSEUNvhi8DNkKwRTwfO9e+
SwiDdSHl2dz00eVIdci7IyAWaRz0urjguUW9K+RAoqIUfzfSNwxaG6dcUwEONWdsqsUaftqHGI5b
aiIdZ7T6nWyA4xHd9ziETHkfP/u8+UhgjRYlJNjXAenoG2NoTUCAY1keCglyPdkbVTFsDVJfARPd
s0ywGwsygrum+FEDsvEyr/95XGftqk53rRsEcB81Bw17I/Co9qIi+ZTbOKNRCh/WcydZk3vkJhfC
8EFd9mukITeTlzw0B6iMyKtaqqoGy3/8HeK4Xh6ip+8yzIpvtHw4Ztljmmae9eRUpHryphl3nqcn
iqL2V3uq66ns4VJGEA7xkTtbfod/i9XnqD/tAcErGQvNoHfnBwJQyMTPGPCXH+0ungu0u8r8gUUv
ln/A4OarXpZquYPBDJPeggX/sAWmDI5mB7ZVFXkxWe464OyZBFMiGlGFIbgMzjdIVomqvPxmLk9E
Nez2c3U0X2Nka37ecCAlJLlMniiaDHCYB0iCBd6qhqHRXYHsLrBOoldIfaHbiJxe538rZHAWfoNO
u0YnUKB9ydVzovaKoAX6LsqsjKfk0qQWS+chC9O0DgJZugkAvdE/eRzehXo85RRXzPhwTVRQmt7n
bKXZV2Sykv7Pr3UMnewsSDFQRaqcrxWycp+QpLJ+x4NdpoMAW9/Jz1N1g5DcYbGZlhe/z7S4nsMz
T163UyZr9nBxZsydGXfn2PlbWyk+lmDwVh56xArwfWR1T/68w32iRd9D8+pgyrDi3Iuayi/YRtjb
NrCTN56hnZEq/zCwEyDBSBck9v4esiE2AqLy2XIZZdocrsEcCLpi8Voy78elzHd0/IMXpmjV9UVe
EY2M9xnUchkI6af1rtztEHmnkEe9gTQJU/zO/jqxkVjvJLY25fNb+v5BaSTIzSD4Yv+gjNG+oNm4
qDQPmhsy9ZPNuEy9W0j82S8n1yKzz9UX1tCV6fRNNVXjqfNf53VcSiDpA7cE8Z/ciXtqEjkcDhU0
IreeXFnqB7UojZRfJQhiDec3/0l5YZxZTu/bR40JcB5ck/8aEyKc+aR6Pj8iZhiGioKyq2Z1wHD4
IolDIMLZP4D/m6QWmr85n2JJkM/oDuodfhP0crp5SGHHVvqawpsRqKhL3LppzQEuSM7BzX8axjjp
ypiQJAS001lXOYjsToUnmLQ0NKixi50HDalAaW0+BWt4pTNew0rffZR4RqB3+XNV3E4bcTt1jJ/d
BAxXDobOXLItzG7rbamZ8drL4/x73/4nXTck/gdakgde3vUYeNlNcqYYrW1lKeTAknSOzzGl17py
5HNrfiVNCO3xPUQMZzf23gJeVJi+2sBW19F8g+uU/bIhoQjn7XBOstCwEMS95ff3YQCOQdD72O/l
h0epkWKgrSsFLJMIdJTKL3iAX5Octh/xWFI5JeDUleNGLrQCRh1evEatcs/Mo/f5JmTfxrYKFv5H
1HAeowEB2CZ9IgtLUgFM8+M40usNMw4nWJiJb83HGdIFlVvVncHYYrxL6h/Tv/aobm/RSULj4oAQ
zNDHESJZXfIDeZ5TgxGwMa+O1OGo0ZHlEHEDEsb7boQ/1V0dTT3+O3SBw5FUfrVjgJ+t+f1hX4th
W7tITkinDt8VHuHDGaUr9kkhInOmFwLOoB/tj3bthw0FXF9qT1WdzuFMwFzcLc+jW56RfoaTJUAR
YibKpS1Z1XwaqLIsNWYnEr9Ieuj0naJBeuRP9sgK44UAU5hkiCEaFsGARLp4PMLEIHOhXvqcvLQb
IyAWlb+DYfaOoTeeFOipllxKisjFv4QvgwWVVMTtaLj5w2mAaPZ1aP3WgaP6c/ji6ACnQii0zz07
euD40sfqO8TaWsk0xO6OAfsW67kLemF/dNhpl1Vglwf91+QNUhOmXDOven7kGk6R5HsjaagBWZxO
ZvSPfdwYTvKWvvyafmAMgnhOV87d/c1KFyzo6eC5mnTkV1Xgomw0EdhYrQ2X4ZcptfTWmwn5d8R+
3dn18Akk14m1G7wpWDjvzNpz2CAaRjdBseEbLVVn2NsM5YlNQ39VSvOBdG6NiXc4rdQJG2kL84+U
i90Wd5eBwkqiBRR7OBlf/21bmmwKFCZqtr7FANUTUCXpMQymPZXWvO2foiztjDcKFAZ/MujrYcv2
45loWTUKvV5T00wzE4nP1/lIRHXcLNTKjVuMTj+HY8K/wh+/x3TvntqjpwmP+qJ2GmHQd+A2fjzW
WjhYIGBIX8L8HJq/yjxGmPh0LZbh4gvgzvjvZhmmT52Q0MjDFiSGtdy+MvhLzt33iYpa2Mmf+ThO
nWj9L8+ZuyzRTAfSS0Bd2qMWJ9bey8/Nnaig9lSgYvooEnx0hZvGcuoNTB517ApLOdKJWVVRSWOM
bOfx6uu0JYX6ANCQgBhu/BrKtkZIrMYZhYLG0ivJebVOxTpl8uDPLw3sipICsy4bue5uakK9zXvj
X6SdK05hbUiO1/MpVyUBHKtb+Yea3LtFWh0v/EJ2n1odnNNtI6Hu1hHfD6oJrwpN0laHjC9PtMdQ
uAzi4qrUSFAJJHyudkfIv9YgBS6FUdWBK48dfr+M1nci9E0shrB974t7+/nJKoSJZXIYe2M2nb0h
6pUtumNnZCNNUn8Z+VeFaGbRACxONhP3y5+jVF2Nz98WU9pHFOv5SPxqnMK5owWY2IGZCm04q4uQ
BX20voMEpAdKbfMhM4Vyl8EM1noT6GRlNhwEzihv94UPQpj9bZAuNTgKS5HqbjOLubKl13JGlxgt
IfTl8bAc1g+EM3IOPzlJJeF5n2QLdTsbukywfJx237Xi9uQbBvWVa6CDdcuE0KrgemgLYcPgZU4b
F6n29pMm4WAJKJnFQjm1zcZQSNnpPg+ny8BWMeSegtu/bBHPG2iZKOiUynkhBxYNOUC5pDC5+3l+
W0M8UEBrJoL+uqFftxpq6H329nZ0gnOb0c5ic/OoUxzJLt7C6VuMGzglbHjYAfIgnWsBDk+r9F6s
35zFDayNIMnMfKDpldk3YlBlRKY1ucjDk93BLN2A3aYbnWfAD1v+06NDoBVsRuiAl69Tu5JfCRPp
/strofGDfnGBkW7SbMrk3sk1EJwg9Nvn6HsBtKxkGTriAk3hFFIMW2tirU8j4TP0FW1LwaoGehd2
6mfUlFVA2Hqq3a1vgTjww/LsFj24NkhTQPknl1BiPV45cOy4KMZtBoOW6M4EQNSMu5Sd8ihoS21r
ULIy4n+zkv7e3MpR/49uKS3z7gb6lA7Ku5DLb40YV9ZpPeWR1cMHOCurpkvrbjTdOIYk0frz/8Dw
pE6ctHbBGHB1lulSRRdfOOVPW1P5I7FhskuFvx8EM2hla9JDmcjgZhtD8fYe88igM9j9wBpTYYo0
GUSVu7i7/yKbh79R8+IV3Kizlp5F0CF894ojs02lwGVQNujiqp4LBq3oYEkL9jSjp/pFEk2PzxT5
dk9cmuARf4VMFUGA4ry78oWuryFzkABovrid5KXTguqXF3PxwnCIZvI5DNqQ0bVbxn5qePwSJ2MA
6oghhUxPwQrcYMM+19Yle8Efa0lTfSWV/FltUXa2tZaGzAdNRQGqKVHuouG6jjaxDm30i+JFffJ1
BhJod2xUoQbX0/VRHz8qYIHMCiWHu21iqQC9ykDwULFBSwmIcw61xgusJQnSPOrv9aJnngi22MNZ
UJENlTuVRzFfRuRrXDrvuYmNonzaiEKLiJQkQ7ej2x+esCyX4wbr7Fy2aEcDa3BtpgVxgifOhikj
9lLkKxxN763Oondz35KfgYQahDMqSyJutGin9skGvAQuik3z+bJbanmRg2GBPBPdSq0uwsg560gQ
dX+5QbCYKvOzIPqAHNOU8j679pgOQs+8tPOZmJKpjAxsQzAA88GImrmpeucElHD3HYxHIdAwMVSq
i8ZW7uqUUrZiOFXbl731wUGTf18ALNng/2fkNerqSWmX7TinKu7/jnGdORvMcg5AQNokHgLeEDET
ZR2AUlsPZJVChxEXO+KZceYFmTAArKx2TuKri3T44IpmfZ+W3//vyMGsbXb1Z+8h0s5l+tcOdx6r
DfC1kEtTtdhBf5LpbuzHtZn/13RW3CcyT44MQ3RydWXaJXnOzpOJuCTya+KEytfvEGqsT6BZ5+Qm
kVlOF58YoMDgJoJac28BQeXpFAa+wUxr9yKefFMnXVsDyXg0cDh3V14TrCt/u67Iy8lHqF8ZITU3
vxG6jVsjn6v1Ij8bMYyzPVlyLKwOHMT1LyauZDYMYAKyArDy/eoT86WV2NDIDZbYFprK0fX9Jj+3
diGgygRj8nl0g81GSOKlG04okAyvWs5beqKlqCn0eA9GIV/ce505eJU/+xfFk2pwKZF9+UX4cKzj
Gib3gEUAtyArHaj5s+eC5avTpFdx3W4FrnwA+OvP9P+wOMdzNuR9jMQ/eC0lrH9Ztu8=
`pragma protect end_protected
