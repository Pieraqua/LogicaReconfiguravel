`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g7XSePYFBidKewaj6FQNWk6dbsdjg/unCWNLjwlpgSHg2tBgpSJN8hu4DYSi7z9C
jxQmIA3Nr++kYIT9Kn0gHizKfvhzn2YcS0bRgNqkIp/hy/H3H6Bfi3eF5Zg43JuL
NF5b/7l6ato5/9tdQbETi23DLuas0KJHvprR7uU4FEaCymUA857yZVerKCGB06J8
y2HcGb0OB96zqUJTfGyd6rVMWdJo8c8EKacLYPa+AttX7SB/QW/XywOSmuGkDvCo
9gSyezFPE/I1orwm/WE9lda0piD2TQVR0UPgNJJ/grff11uFBAHpGmC86uTmTHvH
KfVELvJzxy1BCWMFnJKQOnYdXmmsQc/v1OIBD/gC1W7sOiLLA1qYSCQaLKA+sndd
mbbZhL/+PGGkJlP37f3VNvq0vi125UTb+6cUSVKHG/tcT5FvNNa6SHdAeF4zqQP/
PYE5tELD2s4v1mR6rEYbGXFmWZFaNmob3GmeTqtJ2ADbdM8M16dvMJsUfiGqirr+
X81yGjKPZG8MotUptsLVOzWHRnf6ZkwoDVqq+46aU6mxVskxRIRFRYUlAb0QsWrR
HXUulZBaylsuwxkavaDXpMKF417OO6VpIPxlkViinMS5MmRFF2d01ySZwEDyU+SS
J1FUfuIQxpS2pPLnMvss9zv2i7xGSWyb5t1/km5JknyWjuZoxkematNtCOnzjkcI
7xK1lWguk/l3eBQBlEeHUJ4jASwjU35EMIdHaygEdp3/jR1O69gD754+vIDkjxYa
KXlnfxqYj2tQhrO7mf0l49TT5HcjjpMnC9hlntyG4rmMKE8Ewi21DkHif8nZpcNY
/s5X6+caW1sbsON8ky/zgICxT24yiDwNgAmMo8mFK+Q+mMUiNK6yxzwEoWY4wwOL
jTMDC77U29Xy8don4KM6Zr63CZ/3n+2q2eaezYjYJ3PzGCE1CxrtrpaedwhUfOkw
wdt6IsLW3zxk8lo1lsqWvNyzv6LCyRbgjtEcixFnJ6s77RG56X4u6az5K6uTYEHU
FmM2eZXAnZ2ZTNIwJj+DR/x6kdpUwrvINOnKuXAR8vuKltnmjLgVgWVThM2fDCq6
qv7G94r5rsZX/N0ksi4H6dxYozmPCpDvkYccMmW6EEYhRJRTFBtM39wK9E2Ien4A
8lN2zzKpdsexuNzwASoTHO1YVHRYqlsv0BmuAEUzf/VuzULSR8zd8Jhs5FrWd7Gv
vAh2D+Uw578cIvw3fbxVxFMGZrvyxa0A0uONYK5ERkbtWCF5BqnjSyJxtgyz07am
wSw4pX0ZZ8DgQiaP1UPlKJjL0t4rlVrmEYPxmBMT6f5QlHjyvJswQLeI+D/E2lSW
UsB+lNXHyyD2S00oQ6mlFNqCk0d1qxqO68OD0ZXrsjrjghQ8cY9nZO3A1RrrtyM1
/yzSVyNbIKlHTuKfbYvHMw3hlerqEic1ylcF5/zMgrKFzuFsLfQGHuOZN0w3O0+y
c0MsDbQh88aRWoytmbNA1pwqXcbUb8/qkVuUcpZL9qXyntYVEJPwAvdRXx5+kd8s
+OEsYr7LEciHZb4MwYM0BviYbxHk2dsgsLVKU0ttLQU7abST16zQujIAV1Rn74q+
Kx0RhGoq9akdSGqUjPid+aUiSAUdYMwSx6wCKsOQybYtGefKq68N9X2VD46Wt42U
mFRM+Kd+dM1t8XBAm/FT4JmsszC4olJzyb022rEfs5qKlvSVGhHegZScxupiAlqG
XP4dn9ys3JR9IWNdCfsQkto7QDOlbDKfjSwckj1Hud4OOc87QK0NPCAB6QxjBg8f
O32lI9n7ijn6TtfizUZqjpxBveoak8On5jQf3Oh3/++Zg879Lrmg9RrtxKlglWtq
BsY9iNjAEsDhaGLEYqgH1+/X8gWUDCipEhh6lufYcPgq6jZ3I337hEzci+OcZM5j
CJa36wyFFAaHyAYM7NvC1jLR9Qg+EOWMPBldfbp6n+CH5qFhikiHKo3HYC4lK/X4
pN2IUFJMZMpd77Yu7AbdxDlkfpjJYTGB7AuPFgfXmolGGlu7x7Lq94iYx0u1/zsN
ZZXgRSs+R3baFyPkXP8ORRyoFO3Nim4tBWGl9UEdcuS4gXqcMU6erbxPa8531J7E
980a0z9+Ze0u8Enj1sZ9/HjZUFOrCOO5O6g/xopXdJ0qZtAGJomsH63c++ZF8ijb
FzjyMwAcUIWceZg6QbHatxYm6DdmGYIqJYkioLCXh/bQXkb0OTNLuK0dZtEZBuwq
e+7sM7i2TyV8Xvv/Q6uFgHFfUTBSY60wQz6UvzRsStKnkNXP4omsP88nBiMzyrB9
1fdeUdFphHWVVEiHDa7wJufVMn6fAXkcIJlKtCkMLZy0Heu7S4YVxVIs9yyV2y0D
ITXSDMQW5tasWhG45wSLdJjOvCRUZP/+MasBTVcHrzmgGx8RFcrSyUPqyfRP7bMX
020O2zFuwzOfu0g9awxdgm3iY6lVnpsdEMlb+d9pl//q8oE909rctusPO9yjeZk8
xWR/D71s+Ar8ghFtzZ/WGDQGKuYlnuQrwLUwgWqKRPLFosgz5XbYcYi5BSwBDm3W
qiv/ilR8yh2Qjb9LFw90slwpv3MzjBW9ZsftQKVeodJDW9Dlkp5Sq4vzfF3bJEqb
HICAxt5L/Vk4sRQvGiNAcpDGw/ysgFhiTtKJAozvAXSi18yZnafTiSf0wr721wkG
JvZvGKOhVWkMZAp+kLwDKfQdWxNJcJOWyF7V/xLuFA+i6vPa/ly6LrPMB6Dy44i3
NRjsr9rnPjQz4uVvxbAmYuYsbVNDlofF6fxquSJin9PWN4MVqhSRqeKnCi131usW
K3mSD6aLZtULpzFgsYijUMP7+nPT0oXS2ZEyM3jku8JgC9q6ZCTicqNYjLer1LsA
yVBnMvq18oIUrjVO6kVIxG5j/LaLwffzmLMI3ZVk26LZtFBL5+PT21NDLpJEcxz5
e8zsrH9Wi49AFl5XvBaJ9q2PaITRomizc4V+uimnQ+wbjaXlXnrRS2t4fCKCWVAM
B01cekundzge4qJh3sSlmmm2k15ZuQ5SIcqyKYdriSF3+KVHN94zNOnp/lykg9z0
4NQULTZYPrMShFjFcdtWREaNZN4OUPU/q+QRFaMFs9XnCEZUrbZHJx4wiVUznMaV
60INvxMA/Ob+/L8dmepplzEneI/NuguxBZ1WFLX7S4TKE0pTqYXRYIXGDvQU5wVt
eAbD38elWNoqBYUvj/bUOE8XTOMUkGnysBcyoJPBr3fG1rNO9iwwC6hjl373kbNN
oCc9osk02eWdk/AcEfM8nUDK1ONojKXtQzlFbhlbc0NxiHf+G/eH7Z2cG4CBjUuP
9ILSu3ykprod4CZ8M1bPJMkHJ/qYla5uxa8LoZvKLAj52/XBbc9sQcDY+APlJhXX
E6pwtcVar9k7t0he+Yqm3vMCVxeDG1Ez5GoNlBuRsizfTG+eB0WndeQuHrcBP7H9
Rxfr6ozBsa/8iFLZSYWb6VbqtjbRH5wM5XH2Uzt/mAJO8P5rsbe+t0nt0Df29qGE
ZXsRm+etNYcyGBeFrPPTaau05QjZDjCI5slQa3/BTDhbNtNU5vQThywSWuc7SDG1
SDl3TLmvG60ZguyKnblIl0ncFfwERtFDGfOeJnnx7zr4ZQw/+BX75giQV/bd9fO2
fsUsw4Y3jD+dyuRhEXhIs3SNNbbKrsZn+mZcqghPyN/icF+lwLf7I2CQ8M4gZ/ZX
/PUkxWaimpM09SHDGdk0FUs35E2yw5CtdwT95MscQYPGtBWE2rCBgjHzavmzo3tV
hHipwDfE1pwhk+ZLdaYZlegUbjkxeieHf5hxvK1L0amQUMSbQsn4sxpmQ23KUu9E
DYyEcb7IVcyVUMw6kzIllOhaNmyasZ7NzN3zkVJz87FfXE7N+RNnACSwuZt+LT0I
VqYw3307qwAar9rHIPJMbBTYzIIp0FWXG+EvmcHyThcZqq8uipNJ170OOgXRpA1s
BhtcapkBvX4JEv6Ut+JIFsPGR6tLz2taiWkrg88AdaU0ldO0gEGEAn1uvwBTTi2H
ltYpzDSSeIPdAKoyP3wJQRROJkSh2Ug1SpNtVezQz/7pLEFjV2SYyFSw2NGC/o9Y
rSjNhXrPy0kwOl4FceTwN7F5UMQnfF5cdA56O47xhkFunJlL0UIx6iL3b4V75t2C
Ws4tfIEIQdJBv9B3mtuUKWdsVAXWJYt1sYPWzCmxC4ujoS1EpWCbkkVn7aoa/Nqd
TbfffbyrJ79JvGGvufnHDz/Smg19p7bVIuOU4C/56aw50nifTFc+n4LOdokD+DOV
byUTPd8HvT4J7P+1d8mTGJ/12nnijakFl8bwFTAzWwzcYBaPk5+eFicjkermZQ/A
fc4cRKpB8rDidioSBxUsOw8IeCY0BrL80zXWyOO+qhIIHpyr9rwUTwnKMN4G6/2F
PolYTtjKtIJm6J/UnqEu6M4UV4C2k047jDVoH9fUbbL4yykKl56WogaTk6tbeh/n
4L2QTHKjIZSBFG3qUxwP5dmQr84aNnQjy8vXLRaQXW2ZSL1R1l+XTjjtbquRn7kO
io6WuEaXN3Z6kKrDUNIRUXxWDsnOirEvj8lA7OZppgGBBttgzy/akLW9WFQM0pMY
upp10po5JNp8xeVh5OKoxfrY8CdYnRM6/hul2XH4C15Ce+bLBGjhePBRosLUc2uH
L7UHe66g8ue6xWyc4/I+c6/iKaZVS/NZ3EPZuZ0jQpCqlzpujg+E6ioNDJmtQCOg
Eb50+6PBXFlf6A/4kCGcisONeZfQJUpB8FrPgpUg3BQxHsVTh8o6Upp3MgBEyu7f
4zVU59anl9e0B4qqvLKDgSqMToG8gNyNekAwNGMxTZc7g1qQlMdYaw5NuSoAa/pi
TUuBNKaM7rV5ot6vWdQsBuQQzQlVW4pEGiU7yEdxzJW+xp3Kg9lsU/stvJAGv3ur
ECBJQbQhodj7R12e3L30xrZzoUcuwvEpNq5WDmcr+P3/lvJjmMGH82gnySOz5e6q
MG7fhpc0PEMzJZ5axRUH0IfBkFqYEfOKXsjWc8qJDcSbvlCV3H56d5oeucil75+l
Ty0gXfDUIpoZgd41FvRh9XZZEL+ndPyEotr/lWNjXfEs8pyi6HDLWr7IQsk6E+Z/
aTciwcjGqGeirAjqAgqgwLJj0D20vXAGJmgPu2HpqrIutYkv1AcS577+uIOypaeh
O/uLAZuQl9jElQcIKrx4U9kKfRgU1ZDV+2tOUt362JO/vazizplu8QDp5mkYZtz+
g64x5qsHpdRS/O0qk5o47wiO0W9lJ1B73GIz/WUAEDmh8Ih3Pkw8xx+G4ozFxmF3
CdX0x0N7XONB+dcD+Q4x3ZhtCmhyjVzlBSDua9D9Facyjkl05P8j2pwSv2LSNxM+
a8jf2BQdeXXqKW11xYmv0hXUl0I1EHjTPkdPMKV8mvHbMZNGdHWN7KNq3q6iVC6p
FmOHcpcBFs8O4Xxn7cL2BkXvSRUGxoaa61DOXUI0lN5bOU1ksvo++tDat9hYJQx1
z7vSHXRJeh2LhAQslmmlYAUlwxGMQVLE+w4PwC+dRX0HncVj77QqSFi7qf0daMUF
OFAmtLkpB+VvFMx+Xx1XgMZwxj5ktjR6sltmg4Giw+FReJWX1TJSmsEvwOrnfAAz
zXUUlGNBID2umM5CXW5k5hWREIbFapd20qRKGdU9VGqZvVdgSD68GxR56s89TWOG
32chPmSIvXeJWOfGEHwzkkvlRKEldJG2VTwcQSz9x1SmdpC2epeWATmEIoLMoD0t
+DArriuZ5PZEbazXBpkSnHtkDZ/iuO0nm6qENskx4NxA19AbFiFzJTZr0L321Mj5
hYdQmxQhqVPFJK5jrF7JMAZ5eEengwnUa7lCdUt/RJUNNYzgJCXpwDQwKlsp+AfX
nKPZIRQGa26H8V7l1Gylyhug5xnhecxTiuyZ+dLTtT7pc8+WJFU1P8NRyJY4z4qV
piM4NrnAUv83VhUWML72KImi5P7H5nuuColT5onf3rYN7ejbLK3T0am+mDovO08Y
L1GjF3uX12AdUplm3fOMFqNR8GhoEyU6jtTj+k3WmXKfLrbue6cxhVkctpVVhf8P
n8Ci5NXKdWcMLsqnnexd1zzQbPrHrptVTd/h526WeuIggV9wm3MVYpWM0kbxTqFD
H8aOS2doFA1UR1n2wOkQ1ph6T0+vaCu5aJcsLpLclXZL6cnNlIICHaeaYRh2sNsC
IEeG6HJ0Zq/QAfj4btdAQ4Oian/RYh0X0T+9VXQXYIfSD+prJOCBWDjZjq+DOgYX
ZRwGMp8hdeAquUPe7nnql1uwUJyu1qCRb+sovUMLtrbQgYNI4Q0MUas203wHNGpn
SU+fBvcaSDchv0fjySqR8RXrWca+I6c49Ru+Obxt9pQ9tcSaiLt7IgTmKvi6a7/H
q5wVlYGR28iMrZIVVZE9AaCAQgkRSQaN1DgkwcPDcixi8QaPJSAXk/V7fJWI6kDu
U5pxqr8SstNMRlhIg4N/WpZ/mxAYfNRGdYiHX1GkOFT21yWPwXeK4N7O/Sc9RNZC
eacnPROCI3gEyWfl2vn/1oRFwEaeaOe+1kc7+wxg2wI+xmwfN1wWIE9/YL8fyH4O
ECkmvOZvEDqDSDNPwqM4HcEQSW+ax8i8AHVMifoveb4Kpwo0NQpKXN6OiOZbmQjW
Ge+D6jiZgslokRndl0okEzuhsJLDFzJq0atGaAqgR9fIm4iNlK7ZnEROATgGxvIb
QjLwQ3vcOUCdxtuhy8aXGNaterLR540DQBiRECBLGTDH8uCUgSdjO/kAXwUW07/D
KSHW6vPZ8SYgL4NK1+P7I7MIor2F9LNDOaI8Lf/fIgAZjzwrGfjNfiB8mkNUJusV
TMKLJWu22nJlcQ22pHw83mabIid8eAiMzZv1BnJWQW2K+YhF76cKXFxY2qRp8Png
98w6e5qAFw7gPcMZ7ZgmEFCq4Tcp2upT4xNmwvZ8D1cPSuXOSO/n53tVL6YEeHX6
ryIrYkkcr8Na+bnS2jOJ2w+idy4ha1SkvGuH9Ul3aY2CispOK+A8pGY+GxfYuw3B
4r9TBJ2HNARgGE7OpiB5T7VSyL6dEcdjicK1VDp22P/EQzlPsudEuanE/byPh5rO
zy0iDSjxSphDnEimaW0LYcIpbzVeBq7dGdjT7pY4hUKm1YSkNt9nWu7dGdu80E6i
ztUuVD9zVPUHGEbrCtw9XxTVByitMxk9FL/7RJzIGYU0pCsRQhaAlYpbwbUfPBKC
ux/2EVnkUrIeuMZG9iPa1bAFiiTKrAYLm0hM/KWSdhW5/G2lqDlmv9TTua5W5WzZ
sDrExkjoIuCZ/S7VWpHQLX6kYQCQJvtcjAbOl2euVYjljJ8JqvYUTKsjHstVix3h
HyDvStMYgZAIhHJsQuJyNhdI/BS7vPtQQCfLYEbwTow64N9mrsyQB3M0h6XTOaS+
iCWWqBdMozBiJ1UnlSRlT56Cr67BvoUJrHqhHoCVgoHSTHvj1oswj3e0AIjQzTW/
tMAFm1xVQmphwsQk1NsHeEWrnU1A8OrivUx782cxoZUGyzwIgjpy0CyZWLhmpbLD
+Mz6zuf+sAZUaJjfsGVLXohXGMUooYmA71q7hpCB90Bx1FZgf0rLm/xyvGieEAeR
5vVeEm1m6a7nplIIQ90lPrcJK3ABWqDQ3iJt82bbJDlfJQBNAPPdWUb/gOyrXqX1
/0nOIZOSUV4kxemlVKla9CgHV1XqXYzKo/b3psTTYeouqVrkCihIlxePkcFPcxo3
0U+GqSrDiQ3Y9cmuN2K4H2CR77THT+zDLDmXpTkBYcNcA6UpZjXRldCFIk/xei4A
R1gPmdHfbUCo6HKc5AXFpPLISv5zbhpMZQIvfDKZDykAUWy7C4Y21fNilRTkCeuJ
Qkx7NFyAc43ZufJLzhMETMzK3CZVUwyHjuupjVh0Tkq6nR497L29r8uINkrjMewi
r/CSO/Klid97EBZr5PZhW7eanYHH1Cy+SUZY9rsicWtu4i6MdPH1GkdW14VqNUk0
EBeSWe5QMvhFb90Lxf3VzXDDcJf0aYCpa2OX27U3A3aeo8Lx+lI23oYisnWenDZm
5TeM3GMH9Kz5BeiGGZ9QutcrZhy+zRX4R6+txLx7KGsufBN/mCORZ135LPYucv/K
PxG3c24PY9q8ZFr+mXbXHDI0QFb4F3SYqyoPmttjnbHxwGhokZ9YBcnti/m0fufa
j9e2NzEBk/7OIkEMpf6jPPdjv2WKlejjs+XwMI9Bp/puyiuq5mz5OjUnvsff0bXi
KY03uFmKJbb8DXp4fHa+s5AsGIpb+Iqun6CWQR4t0ctgO2DkeeHUVmFUbBPJKxiY
Fyx5DbzS6KlvgD6or0AwHXyqEVbyDB0G9D7b6kdSKsIXUA1HOiZaBhMzMITPj/OL
sVPzrgmT5woySHHkH281twYwIe7T+lKw6Vs8pPTy+CYYrP42ZUP0YblxijVZwB24
42Z22v1H4a4IU9XgAqwPwI9CPG0tWgrDj4zh3K2LY0a3Q0DPF13fAejjv0noKreZ
Z7gDb9B2ZivMa/Ja6J+/ZR1A60QibRwauBGuJhBv5kFF77y4rktkHk9wqFeeVfxW
oIlaLgFx0Kzq2AtYB/2LhXvWDyecQZBK58mHv+FKSZ+PTZ/BvdjJ1PGLXpEUaqJ+
Q7f7Ocnv8u3gbvN3+xi62Hj11xq7I8FIVIElZcxBLiehHsm24kjbRhH+IOJ3VGzl
d28FhJMf3fvGLm6x2wODQbVFgN2mXqtf9yGLbzi3UDKoFW5O2uQiaCXQEM7mxJIy
ntmjfajSiOeyoUW5K2mpisvImQYMUSP7EXtQpWiUrKClGqrnnxkPGKIdBfibBJ6S
TUlX9+xwZzK5JwJPLjQof/Hz9WauRUdinY24+MoItXfXLm3EXt/jLwtdVV6n5I/X
seJX7XzCfjk+WxX73cazieWfj8IjHZn5PDX+yFM1tkodJny5fSWsUg7vetKQtPX8
KYZbHOyX3YYmlHZ5GiP1TQq1fRXP4DYhK+oBPobfPucxGIeK0wG268EEnWs1eC+C
0vuK5PztXjk5FcbXXB1FvvIRE8JD1JyTQYk4S1ej0P8kn0B4CPTcvO91W3rv1LA9
Br/GJLPKHjnoJV1quqp+Q+LmpdahkOxKqTU56ehsTPj7vnfO8xBlRzwGXi+Typ5L
yMwrfVJBrJv7D6ZFbrsN08vUS0pVvmkzEszoF2mNEPYKpdQVqptpSfwZ2YFyd2xe
C7mAly8VJPRC2k7Q8pFLGTmtp6S+SqQYJVqRxyURM4XWq8G5sbX3AssE+57GtyJ0
+WhMb9EUlUjhPiOr+4IVx0R1e19Ut9jpsz6FjctXLH8wY8LqzCHYOfyf8k9fEKwa
1ggroiUiYd2foFBqDrI37szlEEzURgOYcZ8Ekd7xGGur0LnG8+ukIrup0jYZabIn
FhQ7bHO3hNft0dh9n7wm3+IHw5jSrMDQoiI+q0Jr6ihFpe2vxpUVl+qgHLypviYf
dYO7o+/WK+6plB/hpQ84jlaz1fm5P0x9Z1f5xFcy3NlNbF7El58YmNn9qf5at8WO
N/WIA3nW8qW7thOo0AUlo6fdINEeN8YGlhd1tcEWewJIUWcGMa2iqdA38sDGLO22
p1UKl7rJddJRgVAKIVwlCZ8xwuLUr3A8CUdKHlE5wMXYj3HLPWhwf4FJzqg3b6yM
csjplj58IikbM6syvYVtjYhdMhzkaNHR9ObZ5Bg4KYMj1ToVwl2hiPCDqQ71SRfZ
M2Xm9dGmB4voc8zQDpoTLYcE/oYohuIbEDlnhtqy/wzw6NUfuvV35O4JoMjkioS4
mSrUiJ5tJV90eW8HkXawWJ9Q01FkAxzxXLadrSIPA276L9s72b7yu+dGFsIr/Oek
TrsdBq2mZTZ9KXa9Hh2u9JbUli/sSqqsIKe7K/TOtZMWM8wVCat7X/MTkxi+1Xri
xfu7XBa+P8dfYxhCUhV5YF4PPYEan3ml+ipuSAhMAlgdYSODhBDSxNGy+Dzb5wZX
KRIWLqeZ6/CdyjMaqWuHORbykehAj/egWdTU9zhT9/xU4A6uTX6YJOVDOEHESfo1
mlPTRho9jzDucSiIe3deoTk6htUMeNpfxYs+K5TiZkW6zNNgh42G0LOUf8oRodTx
A6gGViyfeCrBbW3aX4jLjZ1D94q/qgtHA3dHjKrcC6zmQSYAb+31CeqX2YfRIYZo
zu+bScGbmAwJ6lrRPyVjEcV3IY1TIGGmsyWPf+2E90glJDhAJIfKew7+V4JljZLm
KEJdcBBRWON8Ctp6tCjNA1npXDh9jr6BfPa1Gsfes8AT9zW/GIS6r9SFQvLUddN7
owTlWD+xfZ7AP/yBChrjbjdZQ0hJYIvQ/bNeKhahQDSSswhlZrh/av65hi2Gi5S2
lRe7wOy6Nyo0ZxJXTMrBf3sFwL1MbIyMpXqFzP5ZOeVXPBFNxDgBacPG3ONJ6+qZ
+0rFwVyfqDqk6nOiw4sXGdqKU1VAa3IY1gG8tizsWeI=
`protect END_PROTECTED
