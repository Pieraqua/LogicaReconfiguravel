`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r948+O8nEzzhqpLhgCln+yHQrcKJbl8rEGAytfuWJYkh1rIz860dbPU6fO4XEAV7
+DDr55/cdaHgFt6OSb6ScsD7VfWF9wHO8EgILNHaON1rao3EnWNBeLvc1mLKYkk2
QrHhEBZ/g5XY2Dgn/2CjpC2aFuvqRdN1Dyxl3WbFQ6Ry6+HxKHpQ+EHlF5QSX+xu
A0YpvAgBIMzbNz++4gunQeO61rAdI7rJVSY8sjSCrnV+8wCSxaadPuFpLJcXopku
MRN+KYUJvzppap/dI7g3D+317CAAYpEz3IevXt+bAosPc56hYz44bmsOQJeCS2hm
Kv9CeXaA5I8q9MYcY9xq7VJCoT4onO5C9GT8s6HrlfanbZJ1cs97tzJulnTfEbE6
+TxFkXe3P+Gru8bgejbdkI8yJP9/QV8WIRegBPpJbRRVEnEZz7qkCraj+xPa7kYQ
gP6g1RVDPFzZpubY1YIp06axIPzB5ja1lgxZlpQW44y9JyflrYd+mXtMpeipqmjH
gs+w4sZb2G/ZRZPowv5e31Ve2huQ2A0wWp2b6x7NmIAIFgsTkr5boAiOIK+0vTH7
jbN3Mid6qMFcihakWFH4fgV8Gn142306RMo0hWF845u/+AoU9W9gz6e87IRzKpoe
xYsKTl78EE1KuTiRhVYjfica2HIGShibx2eHectcDkU1OxOVc3ehRAhcrVBDF4vA
mIzf7/qFCrRPDAkATBK93v1b0zsZJiALT/R0uqOXLgt9fEPmtuQaLSGOcmozWL/D
HTlUMg2HzlLI/vpRKjG653YXKblNC88ieP1nbkZIWaoobxE1xIyaw88R0BerxM2o
oYt72kCY4HXGSH+D8ZH9CuSmvrRF1HA+wwhhCYl1T2CNv4QtVdY0we3D+0100TU5
1qur5KShYZ5mDX2bJhLRN8uoCDUp/Mh1x8yUhJQWk6UHb9kcwKTfTlPBhrRj/U+2
A6M/dhdoBVkX/3t6d+jjcG8sxKjbocBWaEwf9smm7aou1THDYDMWZLtcWruN/W3N
3oa1XPWgCX86Q5LST8KyhmUclH6v48p6XwKbnru4dFYmbRzEGp0idPFbQ4LS+Ta3
Iig8sAUOmyhNHBsN6+/v3TNLC+yAcB1DQGeHdUfb7W2Br5HzS3PgrnxzovnjgG8d
5h5F1+iB35TYu/zTOXDKRjBwyZ4afCotlOh/qfFqlhPviOdeV1wQrC+HzeSvUipH
SX0ZzJNHnhrtpFE3f44/PnY6ucwl2OnV/OvyXJ1MLh+gpq7lSOrz3p9CNOkYU0zP
+PWf49p14P7MHqCDqKJLGIQeQ3ZKiMIoWV54FhA5/VkivYGXGHsfrpKc9t289WVp
ZbxS0LsQSS+BZN1W+x/tSLjV4LZ8CiC3vuyzvrpdLw/QOd4kOC1gjV+kSYN80QYN
CDZ6hX7A8IFGQWZyseCzwbgz8dhj5F6UrDWmhmGju+lWW7IT3h4VN5hT4EHZCrqn
S4jFtLw3yXsxv2dZkc7M6jI3896JIEEDJMj0DjONqCIgPnszG3YGwacL4WzAuYVe
89unVbbUudTQa8bRDRXwEMiPtL8k9TXB5zSbgmStjZ8tYCCE00wPzAFhKI44d66y
x8R0fwqSQCF4IO11Ww0eudj5VY7A1zEbaV2Vz6nwinlecb1McsfZSP8Ce4Hy8IpR
5KJwf7+7ev2VSUiRlsAFAE5J+W/YTSFY0J0ECUGzHXKdUp/XYra+zeCug38CWhGP
JuANbdjiWAEqlZY4MERtppxZQV8lFXg132foCPnXQptl5xGmrK6KZljAKmND9+l1
Qv24sSden+SfGTnRqNrbn6rIm2NwNG6q04512FnJCTnFY54jou422Ox7jIFUVcEG
W6EPzDyoambGlAvlOZYQQk5YVfx9GDo1Xp62EuVnqyYDP8zlDdjaolA0UDXe+/1o
B48VTYiIqENF5wzKv851L/x2IddDf/J9w2BvSF1xf6ggPo0Oqz8FWNFiwo5BoGm5
oLQQUYLT78ZP+ef7N2UWOityloA4QBEqwfvXLADoc+7sG9dfjc4L7P4cxWpMq89r
AfOpkSxYWnLMOZvd0iiIeDCrkJYXTwjyzd0JS5/7Y3IeH07xMG5Ey5h1Hy7Oa0gW
bSRAN+9GmUgbre3aqriqVvMuMl4HCVF6g73wuRtU+fuxO4JYe7z0XqoSLMD+ICWb
uO3/+SpNtAEfvxeFfId9QuO5Do8LgMTHxRuu+wPKdqMLGXH+ibXRm/XHv7q2CQaP
3D7Bc3gEaCf9Cgfhyq6R2A==
`protect END_PROTECTED
