`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kjb1t6r1xLljHWGv57JTPBGrHlQenpewgYGdCA/lnK8sQQMkNopfopw8N0gfHlBe
q2aV632FLV/wU8eLwzMkwg4ihdtNMMzUnjnfGM5xSkzwmfY66fqrnCfkXXEzgins
ItwR6NBDYaTfsiaONLH2fw67PizCxyA32RZ2i4W0/u+RwUEmAAFIRlH/E4CQKqIW
lkYIxuZnXnEVJHBo2Lnzzy2D4gIIMuEIy3eexFJjZTF58EX+TvIxla5cPsHwl8hh
RmI0FOTY0gryJeIPbMVPz1+vK+TB4GXBa9eXzbnQoRbb/um6JGb9fPE/tvlyRhNq
qCjCzhdG6DKFlycRpGAx4LbEM8bYIeqf6GeltpA/TjHEoE2ZoibS6U2VWEHYK+as
eMgnuXO1pnU6UJgyPp4TVFro/pyUxq2nKjKaWRxFBZ2wQj0IIw4T/nppETKRhtRe
k09TKbl8yHTe1mjBoIS87MAufS1pkeC/43+KtRBAgFGqooZH9RkG38ebNpq9Q7zz
lKax+x9YaquOjgK8mgvqXU/2jgaANJwT5H7e4S3oKFt/EYTWR29Tus7KyiyfpTHg
AaSPDCFTf6O0HJSGplBRcLMUO6Sw/72sRXsvHiQWcWcvAEvb4EWlrGrguQsQun9n
Dc2ssnSmSCVBpBDVM/Gn9i1emYeQQZj2OnwoHwOP3QmXKGsmP1XFC226ISMZ/mnt
QStjzhGgzMTdXRSjaV+IJp7R3W1fHtHBsUheu6tiWPc2nUQQST9E8B1iy20upJlW
IxG56KIoCUYKAby6CXP/4vWjpQvE66leFjZ1cL5TW5up16UGYCZt0PQUU3EVKPEs
FmNrSc8AnAjCrjONBJ767elP99Rx+kGz+sSp1Ql6GmYW1CRlM6qciU9eYVHRM2N6
VO09M6TbZ5rQ+pYm06qArkG8EpO1YR5k4b6RJg7PMC0nqKH0h2F9mCrCxpipv3NT
NyDRn/pHk7VuDJPRifV3up4X20PaaJrNMHyxLYsGl2Slg7ufr+CLV13rOZoqj40a
GtSAh205aNn7m/cFKC46n1r52mEMgBBf4pF1n7qHgIh0nFnAtun1pYJbn5MGEahZ
STmG5lsqou4GkEJvkqkIs/HRyphyd2kJrPTJo7fz/xg360cFuiPUuc9RTyPfGG67
JkDGrPlvzImO79iUA9wecKipmbnua87iGAb3r8a+1fnh5LQhpqRezDXqew/UxnP0
HVnseCier4OS6G4oC1ZvetSSXSP8Tfd9NYljJ/ntsmG6g3ZKSurwWsagMK33u267
kFPo7VF4KbznOul/rptOdNBthZjPI+PzxCXI38aiwK9hgRB0TdCmXch9ShrH1hhs
m4CsWaRCpjEN3KoTralDU7G39CgNA5qN/xvH2bTUEe9jr9BAfcZCV7o27Y8lY4Qp
aidobyeN1wmGwOsJZDsMdTxlX1YjrYD7r8NWHgPSWtccgN72SqogWZvpRgd0wAin
v9pT8ZC7zRx6D9uki3O//o3KFiDGMP2NkEZuJUnmFS+1UYLf4mDGqonkEosqOygi
vStDXitEtYltIu/pHiiHhjU7Skw2Efq+r1cNG7pfppp5P+KbF4jzi35UIyRJIhOM
9R5SU0Mmu8I8s8CI6y8fbDAcja7gIhEfoqhFcD7QTOXEUK3Tn3LxJGqZ+ESuP1FQ
f4YFhUbvbMdV9J4GcLcLdgkJdUxB2Xwm7L2zjUPlY5CLNQKMS3R6EYYkhYpOutMN
y+hYpGw7/bH6M0iVyY4/fqxh23ju9ytLpIXBR4EbqIbjMogWdmCln6oi5q9NGZVh
0rZLV5WsQAfBAzA4H7WURIsKg6J4NtxicRQkPQu1OC9LPsSaTmbdVNGAwX/qRg45
2DKcAaxyScRSlysTUDj9o03x/Z4DqkUPGj1JcfZL4xuCmtblPMDULHJUhQh6pRlh
7igHQtHc9B/YFCwSC6vn1A+ip/fAMGjzi6BO/iB6ktouHc4SRA1DHpedNnGI6fic
sQV7yNkk86zIKVavX7rpjBBN/soJr1FOoX2YZ5x3hZI2AKu9mCqy9LkHZC0bJm/s
`protect END_PROTECTED
