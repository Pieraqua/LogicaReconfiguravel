-- unsaved_tb.vhd

-- Generated using ACDS version 21.1 850

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity unsaved_tb is
end entity unsaved_tb;

architecture rtl of unsaved_tb is
	component unsaved is
		port (
			clk_clk       : in std_logic := 'X'; -- clk
			reset_reset_n : in std_logic := 'X'  -- reset_n
		);
	end component unsaved;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	signal unsaved_inst_clk_bfm_clk_clk       : std_logic; -- unsaved_inst_clk_bfm:clk -> [unsaved_inst:clk_clk, unsaved_inst_reset_bfm:clk]
	signal unsaved_inst_reset_bfm_reset_reset : std_logic; -- unsaved_inst_reset_bfm:reset -> unsaved_inst:reset_reset_n

begin

	unsaved_inst : component unsaved
		port map (
			clk_clk       => unsaved_inst_clk_bfm_clk_clk,       --   clk.clk
			reset_reset_n => unsaved_inst_reset_bfm_reset_reset  -- reset.reset_n
		);

	unsaved_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => unsaved_inst_clk_bfm_clk_clk  -- clk.clk
		);

	unsaved_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => unsaved_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => unsaved_inst_clk_bfm_clk_clk        --   clk.clk
		);

end architecture rtl; -- of unsaved_tb
