`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HJkoaqFxHMiWRPuOtr1YYDpjsP2hUQzlvr52LKM9riuUd76yhSKBgEy699OwH6xJ
X+6MGFpZwZXQfQHpIW5IkLdE62XA8puTd5P2A2KkxNNb0+j/GG1aXD0rFKELBNym
JpHPl98OdMbONlECPMNuN0jTc74ibTfLJLForV4d10PLLjzP96WAVR7tDX6lWEtl
UkNAucMsqTaih4WJJ7KV97zgjfCNsy9xgA1haZSOm0UEE2ggOLP7QnuCdaPVrziT
P+Bfn1Ydaivicxtuba21W7mD5qFk4zeJR2unJ4kBICQyhVafYxCJWOpdPEa7LuIR
GNo4vT8ZXjY7cO6oxLr6hfy7PszVow7YobcCxmJuUzPyBJluvUs0SCHvVeAh8Ng7
b9KOSUsTCscKiZZjEHEg336NQTjKBxwumIGHrcF9pU72K3ZSfdF4uCH/1LXh5xHV
beURpUWgtJvEKGwJK7IbxEdXjHppvxzRHOCMuKE4U3bU9vHnZLuywwClNvT45JX4
lMLO1L8tZZQZNbzTFPC/DaSYLBrtaWdvLee5CbfL6klnpS5mc5wCm/1d6TacZu8r
Y95nOuZvkppVF2SfVEi875hfj99y6T4f+L2G40GH2rhImJ883z9NeXYRxs89TE/D
dyEZpfXkenpqSdDhgRFP8WiYRyQ1jlWfo001bylF2zDQHKfzIosEyqGth+7XZWqr
eXABZfR1CvAeV7dSB8fZV85UaJOMre37+jXiixTz5aZJjM2iKSnBm7+ilbYxjVCH
jOn7ujVceoaQFEqQkMhyBoBEFH4sQKOjs0sViKlNQv4FpRQWQxHUxQFM1AgYvrIw
V+fCxFLGrkLEmCoNmmdzfUaEHwbuWofcwFT7DLTMonyb45I7ONABiqXgrajWt7O3
BPTU3DuN+O0ULiwG+iuwRa6dePynuKaGdAnigiyGoyuuZwsMtZf/P1dV+s7j+oN7
zhpAOSwpHHw9Wi3UvjsQZ/aDQvaYts7nI08ok8YIibNi4MicyQlqUo5uHxb7mwx9
0Ox/+qgJKs7cfLFzFGEA1zkgjwQQDbSHqbSRPTMH9EVwZbaFVSiCXSG00LO1pems
aCUukd2Ey03td19rG/CGYsY0Z9KkhuKU2oQEkmwddn8pybd8zL9Ew9uPQuMhOXlI
2R826eWtUWWkyducxZJLM1qCBZb5tggbNEUa3hTAGH4/hN+Thh2bEWxGLY5EEs49
kqHmTPVV54Co9MBqsO/vxo7gfPoy/Fehz+clwoY7QBwtT+A91FLKkGtbxK2p/LxY
d/be0qzCx8j9xIc39neT7UwbCAgyHYdUES8S8kp+OHO0br9lSiZMvIYauMErsip9
nTaEkNTo0CP3UG0iGKdKxa8WKnh/H51VSe5Zbic7CqNvN3hz66iZ74UNGGN0R8tW
307bUu3UNI4+8eWY3NFBIoMLHmVuZ5EdzL0/maFgsxR2T2up4lbc2IA7BmRhkNev
f4tzdjA/079S5BtMSNmjj8Lr9IjdlAlnok3cjXBWnKOTxlzpb4oHm+pI6MjRBFzM
O6Pt8r1cxi2YEwuoSybvlW7jUXXk5sHyQe9S8nwWoZJ3MGM/pkRfNj/ayb8jgiWl
ocLjCvuojgJ0HDfAUiyJYZOx5rWUpP6dajlHvO2Urd+amvXh9m3T8QlKbkts0H3+
wue7Y+fyXbwCf43wlW63qZSXnXKBxAqEkv8pN+HE9KhP0mp/MWVSN3LJLyMtWnsp
2MEWgRhbk/RBJ0Jox3T7yGlAw3fgJ8hGLCd4+2bHDX4qQSrVEZT8jdmJVCrBavIa
lgSwPzqYCJlB5aW5Pn0YwTqBdu1ZLl/xc3cpfq2XO5HipaGbKDjR04rc0COpkQ9e
tLxOkzFdU8W31E0koO+lEsGCLQO4eWfF+5zchpqe2ylmYOUWBkBWI2zaz0kK5TKe
2PmKqf6yIsOm6Z3QgVHv5Q6+ab12lvYTjIjBkQ/N/WfW2AAd7r8g+jN1We+Xd8x3
BNC6DNEzXMAihD4sAPWO1fzgDX0CQwvt1ZUfFUJmqNpbgoW0wmbigVKuq2qga8zK
SyjQWtbxzfVqjHYGUUK7xlfveHE5EJVU+aKK9vBDOYcYb4Hwx27joce9HMRqtIAY
NZRtVbUFnnT0eCzTZbVRvPGi+0fVc/po25qgOuIlfUkN9Wzcpgt8a+1yAOqAI7Hs
lbHI4pluhq+qJanvePzNPPoMmPDZXIuGAws0ygzLfKECUl6p89Z1YlJ+1JK7v7C7
qMYsdXqHR7ed9w43LsdCVl1hfdUOtdVswDj6jrN2VsGre6O8rHlHBwEz9clqLQfK
glsUEDW2CBksQM6Xnjb3GPi3e9wLLOThto8ipgRr/szjsHXHHXxQMlivvtUASCS9
t7Uz078VzH3SYkMy+HGG3zeLVpYkjjuP/qMxTNKLlx+x5zg3t3Q00FSNbnxz+1o0
wiw1kNUzu4DFIl1s6BCNaPJDNZgZGcKObT+hj1IFx0mUeP9lNJffSVd3V+8Aow9i
pmKrzB+5pqi1+zaN995agGVs9fMJLpq08gQbH9H5pbJJMlXea/vB4xjKsEBd/lOF
L5DiYB1YKUl4P9E2Cr9mNFDWhuNbkRnI1MUFGfjLMN3S46vnMCoYSdJqmWc5Dzz3
FKswcOVyNnUFikvKhGtT9m1Zc8JGgeylXZ+/ARQ+T5klLGo1P2h1jfCGvApOGqOD
lnQsfNcCqdXTjv9Y8ybKRe+VpfpfXRmHbjRVJwxeeTFLyhnzTAUSNzwWBjtEY5aO
v0CLgNroz1OE6Ikc5ZXbj8vK31cCo0VnAOqgJvAQU3dgqXbxOyD3zAIVRGs1GARj
g2x2RJYdFGxS+BRT5DSQpekvO+6QCtuVPf3J3URWnWbuMSUMISFvbX17I8zahKAY
FXavaalV9yqjgMOAmCa5TIm8lZiMi8PjqCI/uqrbnAZu59Gb//kGjM6x7cWQRuIH
veeDNZVzjxxn2Msb/0qhEjQ7j4hluSTO1XX+bLXjku1xr2K32Xg/9fINAUaTgbm0
DxsWRPVbQjK0wRdhT+hhds7m+i2OzQqNnH8JFollV24lkIEKwmMARxVuR7KeS8xh
6TVNHK4qB0W0TTky7kRlccbWB6ztMEkQYMrAmK9nBgZyDlVYU2+O7wEy0rPUWntR
nveBndytPxKngcIDRfAxkvnmLsgTfgaiTMkGTfqNOegV+WO9niKGZyuLzRO1tvVD
p4zI9OSH1qiIJGyg5qgGwCtpwEIm6UpLz29rhQWt5ccA4CLUEF+GjuH0CayD4I5P
xbqkcCDafX3rZ/FBIhS9DO2b8TGyKojkY6OGpdqW1n0707YQDIq1QMWFxqT7+QFM
NPZBRG5vkwMcMda3s1i3PT3JC1BlmeOMQff8ISh2qSMlKe91q0rNjgWNGdJDj2n3
WbOqfrINyBBiBMSOAbuLEhcl8nkNgAho9+US3bCNvtDIpk4gAeYfqP5hCIdnHJhA
67PnN+Q8Lq3NRCOjOM+opv81TKjBmJ2K5kTA6f9Vni7KTA8OFRUlFz6oizcpZZEP
JOf+jzVVDmWdXiXpIquagehPdJ2WXn56GQK05dY7vSFcw2H0o1pl/IwVfcBDOH6R
H5+yLsbqCOgVNiIVHK7MZKJ+L70xYL8rHEMxm0YXFHlfIxVcrr8lhIwZvutl/sC4
zJ689pnH8KM308+aP7PHScKaXtraHRTEdPOX8c8jqR+nLB3R7tW36LhK7eSv3t1s
035Ct6gk1i07u3tKcH7Pbbwv4OliWADmr7CJWfF5Zq50m/hemYrhFDtu+F20NJFV
W1BN2a15HKXOP024qq+tDRwtviiQMPGknnVTOTdZT7n3R3j/Y2546VkKtYIUTmbd
OlJ6pwiXodkj7PWgh3EZvN2gttwQGei35dlKxSiCw8PxiQRr7TTKnbjNb17+O89K
h/zpwLKScI0ln+Kk8VZuAX7nKLmwDVHhiLaT1NZeL85Hf10tmnrdeZ2im7VFHwMv
sjtupze8XTBhwAr2Tsj8A+NgSiAybxrvWPIfTbhT/J1pkHlU0tD6/nLOtlw+GbxM
3T93HuyXMY6ly3DAHWP3DwgB/DAqZ9NVl6ynDb+XTGDS4fCS9K7xeFVQ3B2EIDKS
+cWY7tA0hhjEjZHG+QRwa4aDNNhfEwp0zVQEP7KYaJaQ9jew0n3vG4HXKrXMh2+b
f2bh4Kcv/8DlBzZG3PNNpt876cvfnhudyeH0ushrh1bvY0+jach7TtKLMsWbj8z/
8hloXUqZmxSjtXQKCCnYSHQmfunsncCJcV++wXa8JqCHcRRgGJ12QHaQqbPj1Iac
LJ1JIkU50UWfu9dEMFD9IbciwfR+t8EiYtt34R3sHaeeTo49SbZ55H5UeMGtiyPF
vY/zM5GvoznE0q7EcxR7mDtYe59YNYOqQKQsfIlRD1fOUh/ubPIa2gPLr92u7M2j
/bjrdFXvedenZMZTdiDEwWOY5YmFpZkKZtyqt1rCqg8U3zi4TpN1PqFKHDv+2UBY
ihFM+B496pQto7OSzsIhQIkpa/hRgJDI7eiYGlGNEy8/lu5DOoBbkYQ7LsuE7xFn
kVP22ThdMLL2Ykrq+Hx0h8S5hMg9KMe7E5owExyaTZ2YCibTJwfc0tYvYlei++fO
un7Cq7Yf9BV+a5wbUFlomt9dDUrzIwx7r4VS51uICPeSs0ChQT5Ug0Jq0zahQRaq
VxbOeVoL6El1bDCT7ejhW6hsq+fAFd56ypzz3L+AmWQzWUfoMonuGFy+/vLYVqyJ
g+phPi/auWaxTFk5YD1IUGSk3rXUxxsGUltudOJK4Kzflju750RKBu/B67zBIJIv
be9kGv88/+8TxvKO8YXq/TMdfrThfXf7GP3qBxqo9dDHJ2pJ5bBi2Uj/biaAmyoU
LSxQODkHLAFDC94EPyAWoBm0CtKwHn6f4kxc4Boji4nlrupcwlyVsnISUcjVBWq/
4Ow/uDq4XbSjQOIMyQYvJGp4Y/35CVefM2G///DF/GSfrb8gouZAVqlJ1Vy5LK2R
LbEO1QZpHLMqbutSWDjCtPcAAd7vs12bAvqtPVYZL3Jo1q8AMO6uqBeb1BdseWMx
ZwTzZNpwMJcFwgXyCVAnhsCdHMQ4p1IIodfMV+nMsDdwYXeiuDMVesXDjCAT0n3T
935CGXEW3M7phs+3ihUksrEgjmohk65bxoIruYbHw9jLbPgxxhkklSeMfOWoJrmD
7exXyQwReNeO1LbAWkDPnShYM1PqqzC1MuGiGaDqVxGRMROMWl91b3kVI0Q5hnfC
niPIRWNamnVs/PHhW0mGtOiJOGe9yMytNHJzYAbaN/ZCTZeo/0411PWf3bUbC75c
wA4w6XdYjW8yeu0YWj0t+8g9Mofyh642+NPzABZDhZvWOQnX9AsIhFDudq9OfOw6
JN4MhwqRofYgGkVXhgXnxRy79rbb3LXZ87Xp/9FXbeZqXHkXhac0ZJn4O6eAJBo2
aDJemPxk4O9L+BfwYUr7Um7zQzNumcUWo9OtsOGWvhTFU9Z+OS/L6qF+223JQePv
jgmr1/QyjYsdRJrSuiNaCA4qtCG0dYfChphZgGJgqDCPhvgUBQTquyAnjbhzx2vs
aZnzEeGTWdRm5z8cFZEsNcT3714h/u1lMRcbRiq3SpUKkTCKwjSbtDfu3uiwxd+d
xFSWupi9DGIg57ZaLe3t4z0joSpv6IJPA9ZFNxqpXuIbCFg7CvpqW5EH9V7DrEtp
sxHynkOfx5/Bq6dYftcQsaKG0gnkmjs2Pgsruy5rkq2aIuLXcMSGDmxw7ILjj8Gh
5xDhKxPQv9b9V+JhRi07c0lDGPc01YUfS8oUGJ4Cb4Z4mhxlfx4BBcVFA7BE1jLl
MKFrtO16ui6r6Px2iCwPrhoZKwu+58xBuM11YhKUHL2FBV7EGfv7XpSa/MUn435V
yUR6bHpjSBBdq3vLJQ0Ozm7r+XjbwYZownzNZyDGYgH3jogelzsyNW3F7hzsB50M
bDYrki2xzFhe5UHfhnLxOLJgtNOqJ+nGelb0yC7lRYiZZL56Fr+1RcqdonKTw1bR
i9QJpOJX/OHO/Shog0IGkul/rcFgPJq89SjF+REjfH1tSSz7Vdx3UOYka080M2sY
wfcbfsCsa+VcUFiKf0eG27CA6icJVJ+e7nhU4NwhxHswzrSei+OiC7rVifjfRQJm
03qZeEYyN+HayjBJYmNM+axfmcw3AxQ5zo5Yn6OA0Dwae9YQMTi3y0DogIBlwdld
op4RfjgQyBo96tSQyiC9dLlKtyNiF0qG7km59DPkujfiPzpH2ACJzrUS7W547Rca
3Ezc/FPVjhYFri318CqnBHCtyEbo5Zo0/0fcA8BzH0k3VBVGPQFzSFSuY2QB0QCh
bpbIAwIBN89KomCB2mCo33lyj0hTmwB1F6fkUziuejf5bz0vwu+pXH0o+phntDap
oZJreyRgKNeiykGL9xuOzFI8h4RdkcwzprwE5h8R/xgo+mLa/CNFXKfeZZ5xM5oQ
jKWiwR6s/UIJ7ku34WSta61BaSAupGjlwG+ekHIvowgaz3rexr5rugtNnbL8kmyN
uRfHUevQBOuRt4+4AhTAhwklR6kVdzLSpa1mifvT5/XWl4DJJRJyTd1hYy/beNHq
Mb7LiATjN39gerVMeIuJhio5giNhiLhPywJpnn4W8Jc1jF82DBwZtZZJ17v3kNaC
tl2q4H7afcqU3v2h5RGzXFCGYwIRlNTkBPgptjs+5Jyv4perY770FJsL3dihzQMy
sJdFuaHDtybkYNIg5YVFJYNbxBJjuc/nKJMJBgVkJDv6qjFxZem9FrFlUvTnEjSa
DJffcUwL/urKPjeplaloNBpjlUozgLkBDbaSN2K958KC0Z/F6iWOttDbkzpIGc+U
VpSuFz7E0Qy7cT1lTrnaSRgDkuJK1keIj7xIhxKAm2GCWAP75fZ539YjH43mHWDc
ZwjJ6Wf/Ffe727EVd8QLGQOa7ecDtwrbFVy7Q5I2IpB/V+Rqc2qmGIH6b2ZrZ1vG
l42h8/h6gaCc1eiGfmtEKHfHWNys19Ey9m7PdrjL0rdlNg3PG8DoPSxlnPk4cAlM
O98YZb1hIAetrlQeHAsKbYufGn/59UB1wA+ku420VwsogGk8m8deCcy1SZApAFcI
gbwS3yqysFFDIOKkP9rQRf/nCk4ur7x/mzL1uK+DH/+hzEttn5teTmkSAGNVL/ZV
YPyqirCn0Exn4RiWYWInPuVFPI8G88U5K3VVxdyBdRPh7MuA0BG0jqXBSyTge3+C
of4QoyRObHM9JIZMqzyPzzNvXWlvJJ+DkhZE78UpwFJf8X8uwPmGAsmBlZxOgAt2
5oz8bC5nbHg5gDkhrXgcN1JV1DmNdQBl0P1E/upYknZUBs3h/KHLfX/BUlSAzuQM
oi0tomoNcWcce96LBc0nn/djag+58st2lsGbBSGyInnvLXWhZJI/AhKNy2F76cEB
NyH42OAT4F0d/TOfO3NOikQC7xdrI36U61FtMTFLaE5x2GoeZmIyfktUGywbIusW
pJvK8lMcq317qPyug9C+VkMZzxRj35oCo26ehODAWPC7PNU+oQnRorkda3muMQ+e
Zy3R0PpyeuSfZxQep3UHY0Q8eEIDFzShOp5/L6u6enO+cb2SKpryGtKxclxiaubU
tMEmneD42/xNjFfSjcXFMyNb7vKMPhErEwrTpE4lk19W8aWex21GMwtawzsUpCVY
`protect END_PROTECTED
