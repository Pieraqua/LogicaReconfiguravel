`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
n2h5Wezi+cNJ4csMwepjgJSH6unONG/7NUA3aVcHj63uepG3yJETB9DZ+KLOuzRe
mFBZLKhGJhtHeg9+vXUZkFpWUFuiUx1xAJY91AHYhW4qRjWpaKNGMEZ0hPz4LlqK
ltiHsT6RMnzgWjCt6Ptvg/FXCj5wbEMo5UAXi11CUgY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12784)
inEBcxFOyCGV9G4y9A/t8sbQ4b+oJVUSXrnf7v9WrJ3eTKylXBGvj9zTeCuX7E1Z
8E5ee5oxeK1I6QVlw9X7zM3ENgOe6nj8MkiQ8jWQsOG1QS+QLwwWJQGjVPgABRSJ
lWo17u3Cux9bIG2gGc4tUyVofmlQU6lKpWiz7JsgqXgYbl35jhvNjVkskoorzUUR
dLbDX2SVtslzYFAEmjeXFPm2xRJwez7Gr3Ws4sD9XL5wpRoHFEiq/TfCDblqmNRV
pm3sAULiolLhaXpX4sr+lF0+CMYgEsQ/skXqMZIcj/MonIEF1kg/Kn7zEAt0mnBd
cqPjgZYF7Nzs0kHm+St0eRE5XZJnzgZF1NMHAV2YhIb8eW1huqk2SEIJIimmWMyB
gbeICBH0r4SZEQvdsXWOpVrfxlq+xPGCXXV2Spm9ZYIBR64zjWw7N1fOak3B2ZqA
wQXNggiDFoOGTpBvfO6teh+DG94LbsSlrEtMepBE53rOZrISfVzxPOEk0TDfU/+H
kYRmAKOhl4h0HOtNpIQlJv7OUCJJpsfhFma+OjZu4509hF6jbSMXKH8mwmh4Xa32
uOPoJOu06el9VoMVpv21XF2CjqbumIgYMicWJZlW8/6pO5H5HEVoy0ElsDz1TRKT
0vDKeyUwr1al3+S/0kCyZl7uONEy5q+5PJM92E+7e1wIez+8rQAdyy0op1FaBhmN
J4K0Uvfd7/54rwxn01wguFGBUbYY6TouC4GHu1tkCAwDoFHFyPrme95gyGkfsqx9
nrLYXUI4nb7EeVuGDphcUn5snEBy9bTYceDnM6b3L4nRZc3yVnN26EnBISKA+1jN
TymY5IzyPHXGEEN8nT1ff5JDFHz5f8gp98doyeszfkLjnBfcoGk2vI0p5KTiw7+m
YEWtsARr3GO3+pXKh4b4uS7JwrtXcjBk7MQ8eyg1bnV9jmfYRvYc/Zil12LDHjD1
ewtSWeJ/n/RZc6qtt/IgypGMDVKFK6qZtk5ZxyNPPo85PCXN5jscrkdY6Sk8m/PY
zo4fOyqrhp/DEQEdwVyEZANY/+wNUphRX020viF9CF5B6REdLGmHkQN+3DfbyyNn
CJVeqwXl9dtKinzbiz30TPL01gZk8JpfnZs8MaRHvcCSYuYu8GTtMN09+SvTpL1x
SydwB/S/5UWEWHCYF2xF08buVcgc0/+78tSRzJDM+/KVF45+rbxhckwB3ZimKLQk
ba0bUooLAk6KNf+0WHXNKJ+BXfuRLKQBvYPrxde9PFR8NN5xY9racbXXLhh5ieaz
F1ItYgjWVBjh6qVEj4VAg1Mzonz/jPwj5y+3oA9Z3vPUXpPQI1LUtcsNKfTn3hnU
C/7ejwHu0XcLEXhlWwChwLan7VuWXpL+MyZLckthWkXIOUw2vaU8sy/hDj+Tu34Z
OaBtDy86LAJIqTBPJIPhw5Yfz9dbkeZ1JmF0ZziogXZaYLL9FYxg6rp5nYZ6W7/B
ILPKZojDvrrmlxUOnp6bx+rye6K/l9cs8UJHHC0OvWH/cRrXHms+gSTZhvSl3pbd
ZEWBXE0kDAhGypHV6dI0h3CipNxbkUyrBkAKCM6zWxdWmWhI7SENe71I2SWOTYeR
ec2YxUQI4cb6USsdQHG5CgCoKZQWzz5LVs2aDktgoDaN7Ohj6iI2U7zgSa8hLSoD
9k3trN82U2gnBRvFCBi0ULLfxiVfoj+eh5xtZHdNlqJHkZ8yJC+o3IdPRDQAOWsC
fvRjZtFc2CRrIobhcD/Yp3AA+ldxhTIirikClnpEyChkjoeuS1UTi6PyTvM6HDdz
+H31xwCNivNGVP47rzCa9DRnyVr/97+6ecvvIyl1TG9t9QiCUPIwgBPJXXTXqBK0
yGDnCKVrWCqd8C9qGJFgROSyxVr/q0QhApKJKZ/vIkXoH2WtZ6D4gCnGMqZModwN
m4ATuBcCPGjL9kaFhmbnhqc7hHjriWOnFt5oX5HfzOU0615Ct93xP8T+02mCrQ7t
5t3PZs9deLhYBTtxOokio+do42R8NznQWErfRFoCFo4VBSm64CV/+OPrc/mIF586
omwHLbnFrVbMx0VhaCtfHnqsoKF4GnwYk8SGsgrfR+HA0ynSTRd8Wrvg/UV+jP5Q
8IumLzOe5lVxR0mo7Pi2Vcss7UhEWCA7QnpnsI9rMtx5cc+dH1l1q3DgOgEPuk7K
g3B7AbEfVi3q1zR6HDx5x8Ql6b5dCNzrYD9R0I2zd0vCT+igHSni/RYDnMmWGTXB
5Zr1fsnWXP0dYdQpvqNuCoGkqZl+0lzIGIkmUHDCCqK5JKD7+zqqFWQlv0Coqg/5
vCkHb+eRB6G/91aw1oavHHG9Lz2lUrn52TjUCvvhY3iI9Bl56jh/yvH91AIpxZVP
VMrEFQPocDCzErGu5VJNFdnaJ2QXYA7eSmLmmeJl/ECTKFi1ezslTWCB+EG0InQj
xUjW/wWRGl0N8ljKEuTiN4r4depCR9MiE9TN//1RR0CnN3wqSBUGph0A6k6N7LYY
4I0WP6/0EkTqRRN5BO6QC62pVrY3sWt5wb0Ed7EGoF7joCGvqpjpc2dNBHGLkCej
xuM5K05nCeAmUmFlMqlkOQQyJw0K5ulYzN7VfXw+LfhAdyMuYxqTC0pinxRvv5Sb
VfJq/NOUHBY0NLbzBeHFOP1kGBejFQUG/YsD4PciIpfb4sG84rkhBj6WoJT33cbF
dquSMVAeg1TIfFJ/fnDJUFrVCe9COKvkLtc/2ntxvvaNAfvIn4y00RIPXL4PhaZ6
oM6jq//aEWVlBXCmSP9SbSjIrY/ijZ5+b2u6mYPYOZrv2rE3OvJN1sclbZ+zTCBm
X+5RM+NtCUq/Yt8huFRkWuPp+dTYOFKX5th0kzjpspOr4enL98jSXmyPNyE8Dzkm
WKllloXlMHSHB+EOto3Lx3vaw7nx4Ou4/xVTYhjjtTi6q5GDVCEUXg/XTaF5veNn
cEKy9yEFQXO2CHzsx4T/fpYCm4YzgA0TLp/YCYypK8S2crb9HbBGjm0s1So4nFw2
baak42Qs+DokUrVFCnWIYs16mVLhd2UUxMq0SeA4j924kbV37WHEwvvV13piuetu
xpXn7qaKr2/uzwAepOt0mGJS2aPvl8FmcoOKCLIFnhIi7BVvnrpYx6EVP9pRcR9p
NzPY3ljP8/wgvBOQs20qe7SwsRyQTBki3fEMGPgTen2HCHCTjEe24AiZAmrOFDM9
jsL+FTNY9RkoHKAWUpiWI671It20KuvCJnNQb0JGBeC+H5fII/+uVQMYF4Puaq2P
cm1GXucyTghQFno5eUB9se6nqeVzJRoTwwoLv8UgfHVCXJQJOAEsYb1O7YGN2uyv
cgIqOoW928EK22tTaHp3IT8Nxx/wvSEuu0QFZARkw/tTlUhH1aysRAj18w9VDy/d
C5kBQWp5e1n4r7OcIoh7KKC5wp0CPZDceZGu/3gi3nMXIZcsMs30jn4LIV997irN
wTWir2XHzngF6sQlxxnAxbyMYqP2//2bJgCMYw1sCpExim66Fymz8RY+kuFiF442
yZ4+BYTyId2VmJ5+l3Zrb5euE5bycEP4mWKZ/faPNUBVQVz3DImj3E+MhGqVGLBi
EpDHIr36ugzOXdr8jGjbnUIYuBVSbzQdcF9ai5PCRkGYIcT0yg/lD5p+eqBjyyoY
+2Bbk9SAFCzsi6P0HkLEXsyIOMv+PEf/TgJc7CKMPMbTndHo2RWPKV1uYHHkQ7zm
1U2jtwvxsxslZTOm5UY0y/+yxgQ6Hvm57Wwzep6nW2uFR6Q+i9Hz7lcnqE+fGt/F
NAM3DJrgK3QeVkPaGBOwQ7Wh7Gcdi8TB7Vl7hLGZbv9nDAoloThrdWO9UKBo1/67
ZTMUIlzCKAzjoGbYTs/0ZyvypJ9V5N/9dmkBzwcGuHVjDEUtg+t3fjXeeVAC2wF0
zpLHV8xygEuUBsqUievFkZZD6ytSbX8jrVLx6IfmZJqX0ddwo8LjmtdhMP/uD/st
E8d6iAcQzSYkLEnVyVK7f/PdRYvW0NFWAc4AXNBm24R6lvaNvglv/3oFYOCZjHTz
OxgQ/gcmHUMCYjF7EV4mCV6T0MQu44DF62tbsrV4wbwpiawDQl0/xT7BhaNji/RY
tTdWRwtaXVmNilTs+jYO5d4mXhSa8cBkoGugRYSp5lPv/LfRsMlFXqjUtZzWb99H
uPGhH43ERvf4irJCVQZm6/+0ZSwK5yYGKxJQxEo5WH/X8+tpNef+UPTS8rVgJS5O
726vcDDRZCi13gt6hWNDojGivoJFR4iq+U8ID5frNvke5v+Ix7jAL916sc8vz/gy
sVQ/x0w3tTFUNquWf24x2F+jGJ/RFJdqI7a+yaARTtEfwctDvhT5ObR18ZeJABD6
g1edjWAdwuhy2Cj0GXV0PbFRjEaVuEuThjMsLp8jTE5i5agCAECCF9/ozzhBwxoa
bEUdtTpDOyU8YBKqegg7KDjbYQa4ItU1io00ZAYaqdnUO5o0pxhJeMGzgDfQI4XW
pykhG93Uugv74pRnwcEjju9r1szIJLa/C8fPhYRq0CE5hAwGE80KpkZH8cmrXHb5
KPGIxNH1q/MhuFyCzFXtCSFS+Og5M/sL9u+Rif79Nj8GNIQak11iFp5ML6g98iql
N7WKFtb/7c0FQaRPszkxcEwPetLwdntLNdGW9QWfzY9o59yfs+1S6jHSkgnIixub
l+04TMnDTJe7LBF1xl2UW8lt8p2sAtpJMdasCh1/rYO62FvP9XYnfk//4usPs5Tz
GoZX9c+6WFtpZra5d5FQghyqkYSz3U3uQoiG7Gf9gk9UdN7+wkTWwaDFM2Xrbhyo
Dv8hW8OtAEs449BOtsjl8U70llVcV4iMUADNNcc4Yv76NQwtebDxRBqqfv4WiUSC
+JGXVidMhg+efzfNn5KsRJipM32O0Z20TNGqttLeeI7V6E5orWUMB0EHpw26bKZg
UTP2Q1j8W1hUxmDMMxob09qQsdBCRU1jIckLbIqshqV1HawikvKappCKVccJU5Hv
dDketx1kzk7Yn+bGqMqHh5ul/98somK64Y3Q+kCspSO8C0k0k/MsLxXOiOn/+sV5
YhM7Tbko6CKADjiEMAImFZ2LV6x7kylwjwElM5FUW5ypNNMEHxXUV/CQKfodg8uJ
0dDSLi67romXlGXVDQ6XDE+lJBJA0OYjvnOSx6lg9MpTlP7HcKcJuv+GyylQZol7
bN5drcfvqOjpWcQkikGXsFI66FP88wlF87M8bmf1awtJlTmOp4S/RfiB6iFu9YvG
G2UAwuNv/DWsfVTM+OfEKp6/VH2b89tjV6OP2favTFuIYxpfPsK16mLFgSLzhqgz
IgUG8WdE/OxwPENY3VFRU370M6Oba53bo3aoS01VFwdmkFzejklDM0M2OIYDGx7q
RlgHAkesAZmb9XWyCwqAdkRVFeJfQ4QgwZZWOZlQVUXToxj0oOxQOjOeiraHLfHU
HfovDmy8yqDqwoCuCwEjdSnl4FHQtNbSZ/9xzbR/LIlEvaWSkfShiDEXi3pMprlr
2eeF/8dX/OjuDKp0s/kvEQzhAdI8HZgfx7KbEARsEyF1ZdVmHeIy6i87RtQbZsFl
dlYiOFl55OlRt6t2WFsp7kg9S5AUR6DHVAJxKOhRJMDeUE9XJ4tvvrLVPD1QPRBr
xSYAoxr60lx6heQ1HTakU8qll1/4yjc0ySwkl2sbpxe/LS2GBG/Jts7jZwdARqZM
5QvOBgyWFBfsLNpIPhZnswYxQx+BSvNwi6Nu5hcJVeXqE3SWpXM6tCbGyGzwCcH6
R4XbqCM69B0G18n9WJewSsng9MEYvbmLku9GO6QcyC6qgeyy5rxnmH9m9eWxvbry
JXrkqbQNVkIec3k4+At1BZ6Wo6foRzW+TtrmTJ0Q75XugyiYK2qn7RFfLFVUQ/R+
xHiZeQFlpltCcQrxYT0BQA3xhTx4Ic2URLMUxidIXRt7Arq7QcGE95PQ4lezH5HR
VepI61ALaTg/WUj2R1GKo249editOXixCDm/VeuH3EyVNhpcUArdbG00lm+vnsZN
r8rlSeYrau5ODDRcyYbprSbCU5pvoOJ7l+lgUc31Gf177K4nafq5LHXu0lD9+2qO
V7E2GVGYsILC5c8qHXkTbU62a6Yw5BLgscnl85U0MlOd/B8t3RsGL7a6kXaVny3X
qzYFETGQdaLAQBDqJDm3atcC0jgugHFzcXmkRmmtQ/wYt49n+znwmeJVuBjWPcPT
xD2AWI6a2zzAreroFg8oGeulNicUcWTcndWKSbhhUveShKeP6aKni3g4QxfBfUd+
/yqtvbgWvM6QyTYluvwGysLy4bnwCBWvqM/rXAvyLy7qTgcQhC9hoxVrcznEVTjD
/uvnKlyWhdrD2OkTEQtA/3xdCN/OUFmOGX5qVERVsvPXTZZA96bONTsWloggNSzG
cbCsb4uBeUrfF0fTCZn+fuci/AWtcIvDmwvAEyY9OVG55CUVGKimT3Jg4Ky1uaA9
uuJshnlU/L0118mY9CJfFm+oBo6To7iOYQEZaGvBAVeIJeNJ7idWIBhBLlp7YqGw
YrJNGvERgkxYL8Y16+jZVLKwlxy4wGG77zHnyF08WA5th9+tEPHBGuvzVe/X6PD6
JQCr1iAj2iKXIYnREsn+J7FYvD1ODg2EsW9Zu51a72/1nDusHGZxV1mHst/koGHn
1e3LzG+Xy1NJcoLUrKnk4+rqpxu1/FSs4CoxdfPse03K/OIvs8tZGuDqmab5yEyo
ItNi0cKAg0woHubDSMQa0XyAcz4fBtstLnH+gmN+tFqHa+5OErsveq6B9zsLJ7US
O+JO7XumzbJxEaHmU76k2YLdgn9T+mN2plg/qFMh7fee9O21QXwC76ursLHoBAhc
uLVKcEUnpjzog0nXGBVg/nuuZuaVUzrJ067Ttnj8fu3r6C856zPCCDYrtqk7rEW3
ofRco8xL4FoNNuF7Uijo8+XdIuSqHaSRPXmxgmd7tCVNng+gn2fuEzg9t0SHuntZ
3SGKGVJXYmo1of+ru1R6vmOqHM3mUVk/2rp23CzTtg1l8N1YLpvd4To9r/fr4NLH
SyQLre1oAYFAeXUlSEM7SwIe5+ggxXTOdbHMLQRxjzyIoUJNC4/FT98x1WD/rRV5
ILAf/j6QOGpth0YsqY3OgP4aiY8jxRb/ZwEUm0V0yQqBhTiVxL/PqBw9Q0/fJNfi
rLmGa/xLzxBjVq4MhRifMAD3sLWmKOTEocLUFO3Ujc+X7Kxlsi4vo06TkiYAwjyY
WpooIRDWmmiB32nQqQbOb1P89mdlAFueaJc9SkVtvnrXlmRTOX1X5TdnWNnbcs5Z
098WMeCl1NlTn5bH17WkhyM1lpfaOFYYgJVE2VLgWmdRL6Cfs1D8eHOLbsVSP2vz
JuLC8j6biRsLS5y7fR+N5P0EIA7vNZPnla4P8AfM4SVm5EsTgXlyVy3h+6GeVYZR
mpr/8AbgPdblALT0i9junwTVWRP3FTN+FJwDmnpVpeR3Gn2PJW8RVb32F+ulejjH
oEihDmne9qJfnkDuokJhNkZUS6QQ9wpolg5i+xTHxRNYeYeXWNdqeYXKk/npP2Fh
pBjiGA5YEmbiqhbteusc9LVT8AwXWUQkQw4DdwyeqSU4gdEy4U27OVmrrAyHutl3
FUBLr/YG8w6Dq/WZKXChbQkWbMJXxeWv8zhmoQr1juz2PEcZeTvX2HDUHAXwZe8l
6CfQGWWRH8y8Ayf+ZWHQh0FvfQAN7qBO+Kr4Y49V7oMuvyU/dPTiEj2vpj6Ngcrf
lW0I02VwIVb8IwWUnita0bnirLgMmjXo/vqGtl96sGZbGDT/L2BjErXQWzWORSB6
WPP4RKMm1Ntn58i9o849MDUdSR9hk1QMVwktMk0ouByoDNFV2VrZZa7GRgRopbzl
/CsHSaMxm/1dNWOQRzGerQtorJuUq637C3SGTF1/jfF+lPKvhHTlC6WpE/feSooM
LBv22k+FfmSvNH2vLJAr9uOadPE9OPDd4xnKbsBq91pa3YR24K3GQRXvJnaQK4b9
+Eovu9QxRH+vv1kRvNlvqGqYFojNicSjSm+5JFJvq28hWBK4sJw51VzgWdew28W9
HvSPEemA/dysRS6ik75WEF7NVxIzAXfMwZTr73vJvZSPhxxp6EHX/L7oOKm/GMYm
/BbURQaVacn+Hq49Dv2b0hDFh0RKUdoj7GfFru/5pwcAfJcq6rfc2xmFpx1u0GnJ
zZkWqQ664rWjTQVZzKljuossSEH77eBim+IXoMfsxHKEYXM9zVbIZU5McTFxMOVM
ZQs3ndDgAnp5KkhvGYroTYwRTtJFMnTb3+KPLrx7IyNnOWKGSjkxN1wpnpy/BV/V
lfKBHoIXXUqppl+WrJOYLM1ZAZYy7N5AOUwdIMDNE8c5ZYci+Euf8s4FTFH0xzlf
nnO9ZltjZfUYostfWsUJigAIhYlDbbr1S/4EjgN7wYYX/WF5sWZJESuaQZZwiCAH
MbXFaPJjT3YEJiiyeN2ZpNFKo9j+8F/MezRSHy1hi3vSdO+fXOxiFQi4mjKRtnnb
7HJIRe2ux4foxkjHB4LKgR2d2BA3tSZLuyAtIpNgHRPjS1mqBKEs7piKlmiOU4vU
6NQ4WNCh8Nhh6K5iC/UcowqnHA+Leg0ivp29tNdLjDhUxDAZWDiJ7WhYnbOCBTBk
/2MuHfbFRbtWq7IxSVeQSoaYUMoQjm2C+WCWqHpqBCZVT64Gtov/u6R4OjI8ZaUa
0FUpdOZI1ngDHXNX/xSH59wcOvwrTzzlJJmoTELjFIll8stOFL6N2g8mbKjvbiWN
eIE8eW9FaJaVLCZHoz6q1Kb1J/+icGr5PrREeU1H6jz666y95XjeWFIUY0OoCvll
ln31tC7buKZooeCv4rXxL7HFqSA8QeS6b7wYeMlOTHr/4qYdbs18EFCGPCcQbWKu
XF3KBhkfqXb4LQKKH23ii+LSx28fyiQdqV2QflzywRsIBLn9xgxpC99DPZ+l4Fgd
gsYKyALlTnucFLkpdg2x+snOZoQ2NzR1Rmxa/OFz2UwTjZ6fMnOOFYGIjRJyKyTv
y83dNHTp8EKpNngHTmxrwV+qzjU9s4gsBuRrS1V8sWvpUfhe3aMDHfAsSHs/RGnL
dT8L6lhrnSNN1gadvW6gh//2dH3tZTTzP9CPUjGCsHfSk5V/Yi4zH+3BKAPpa2Qb
hIU003tdaiPLqiCe+F4PB6QHChGLnzoUDk3Fi2xL+MBQUrog//6u0lVJrYnMdigY
mXPKDajZ2N3q/8lihFoEmmtSCEhftogskcPSI8etMHTmrgQxcWJXyiBeAZUBpNOt
VSEG35nDf0LE0rXjh94ph80VXD00Jl9RZGcBGemkFcf1CqRIV6usAX8Dz74Lvd2h
2J9NY6Hg+9ThHOsdJv2G9Obao0XnUCsvvgmmz26lbA9F36doiC0c/3qhIG79Abl7
YPpX4ly4cCiLkHNvg818c9V1C+/4soVhV+g5/sMuhO9y++0M+4ISNB0fAwmJrJl7
JdGz3liAY8ljdmYZsnI66SvwlKbMolOHKLEW2W2PYWD73F0MPo/7pFYeDS8OlQEY
5l64U8YHOm/R5S2+AteO0vOSN16Qky3utr39bvy3jb54Qc0ArfrvSbXyDGiZHc45
HYsTDBB4Ct4vdYtMPotwokZT2RHYlQayu7QwcVGdZUOFNL6474rK9gf059h+I1ww
Wfz8dG1Qi4vElwTg828qlirLp05q2ipJ/hsA6CrZl31jGyxZB7UOaKgJkonulSDF
2AVyA5dC3IVn9H9/LkksBuIn5CuItCw4AvYap5kotLx8awhmxn7TVc1eZHn8wyDh
4CS1SS07jN6AkztwwpDyrPmeBxoGbZVPqy09ps/HG8p8P3RGGi1odKOxVfr/D4fF
7uF5jUtbBPH4zxwUc17g/NMlHtP/3+K4UaJ68DFYF1GCvAvQ2C5HpUHkuN/rlitp
EvRkfz8NfCzzYic+7sVi+ZXVJGMOP+WcsiysFt5DFz9l5LTM+4/ERYuAcMK1giEj
gwQVAej97Zhodp70On2cU4XOoZ1HXNluscl+MqPU29k3Hf2z5MrNIIxHg2768J+w
Lrn1JRdT+1Vn6BxFt8kYAVsUaTeNr48CRuUlmWE7Aoh2mWz+DK56kEr99y4pLHDR
+io3KNLWYubWeD+A7Ls9ORzWFyHEbhpKhk6giQC4gHXE9/t+GSqrh00xlvUSDsgG
aihH32Sc/BI6WvlrWLvln3R1Khg1wlXRtrFc0jcBrl+mPzZksRegQh0iDPmRDoVF
ZomhzSOakEUddGuht7ES2ynIoasqp+BitTrRv3gF8k9ApPmeeHbX/QJK7tnXDQ0/
QsrqDE8fXUIomHtRR5UREYHzjW5kq7sfnmBsNkH7OBEIgKqpMMhkCRw4d8a6yzvx
WjQccqBZti7+4UQj3Wo3/vA96vkxuRV7kWO0c7H7yJXYERGtoGLiU6+vl5TZoE1R
zg1TDR9aolMdS98jcIiIElvo3eTTW2LGvPqPisUG+NXq8D6ck499qG34DH0zQffe
ZYEWABm5kVzmra9LtK1OzUz6wJjfqqEU4dnr94fvLeggvesAnNEpSeoCOvPIe0hB
5HYZtM3Vgb8xrqYCb/7heL8bDSDb+7r8NkN3tyrbQNOxpYv98Uqp1gF24PrCx15M
hpJ/c0op1hSL7wOFbxW6R7Gow+f9lnz6YDSKuI6BmQ5OeY102hlftTZ6/rApqlkx
lzdbbbCPRgTkAZKWFDUogEovsQw31coxZT5HTc6CGr8tFsdLWIxcsWpIAX6z5CNl
6qp77IKPsw0JZajHCWEUKoMIpvPjou5yz8SMAFmVQYFJ4Gc1itxXuPM1zg/ag7pv
X2lPdf5LWd5PDW2lWzsqBMxkwolPIF/QjKqTBJrbAvL/nD2VlkO5uo68ofL7NHOS
d1jRw9JEalbNXI2/WUmMKF+1cs/UkY8DifChLsRtgry2r5TsD23rQlnN7ZeoAJ2h
nm1YhBFaD85TetypAjnR8FL1egBUSs0k4MNJh4erVmOqH+jy9NUFzfi0TqXivkq7
QudaVw9TCVYmq7t0jSLQO7gHvoR45j5ECSzq3d+Vi1ySB8QukzWBw6kb0bFdnK6k
892hArcAKP5NhIN2V1JvLIDt+99zaBTecsk2+0J/j7mqFuEngLt6orCaIHKQI02y
OzWUbaY208rF60wyhHytEzcFFANZueDCiq5fk2/PG2hXBA1kl8Wb1Nd4h8R67tbX
16ZaDg+fEaCu6drthG30gN2vV6ab0YGvAqOfW6VzY9ZvYmQOwLVf6WHzaGpVIf6Z
ha4IFdH1ow4hN+ITL+xbXYRyB92EE0TI0lJ6E4AUXASeufzfc2ThwVVxeeNvr4la
yeiyzIObFbpLNp+goU5oeGkFXM8aEyOuhWkhvIi5sRp7fldz7WV73iZxy/hvJfWl
LgnRBWr1XEVcS9M27y9hEuiyCBj/ndhXqrm7dZ1/3a5i1h11NFPGeBD7ovVF8FKB
2/+TW+Oe2OdJ7O7Rx5UjCN5XKWcJ1lVdTIOc5pI4hjW0qRp0lx7W4eJ0+4F4iXFM
knKB49hGKa3o++UbVmKScwqPdNUXKg9N8385ZvRbiRU/9Z/OQOSLdWB/qCZj22Ka
uBA9D0NIoKXSxVXQPC0AYkOtTEbXB960J5LVZI8YB9FGeQYxEi04L1e+z2dRJjIR
1sf5ru3oGLJGOSxL4E+cLqwsGPp0dudCdiaJwB/JpJueGmmHUJ+HR+lUwbqp+tol
v5dFHoe2Vwvv30lgHh56GvU+q7xh0JDJlPai+nY5YcvtDgOaad8pU3pN5wfx2NI5
7SRLP4n+fVxbyD5F1BcQFtRcOQHilRmj5z15CO9N4pq/2livBY39bb4X5vCaTAui
EG+Aqz8h+5G01lqgPQUgeXKkpPxUU4RY8mo4CLIvmMlXUdSAZsKDl2uGuZZh5+dr
FGIqjCyxRlV34STYWilVzgCf+ZZFMABfGibHNPsOQi+Unim4dim/3NVeMmeUSuVT
DuEyskA3GI6Mf4k9xpBJGXPoB0FbPTKVyKyhXjScNlBU5cWT0zKS9mmGcmZ/w1qq
TXWuqm2bWnr8ku7vubA+zy0YAaqMQr5Wxv7KjrQUKeKUP738dkGnim5a2NeE1JWG
h7wPs9IP2Z5P6/HrzgG2DiwXQaqshZrVX0OeRDgpBigrH6/j1B3DMXMx03tE0rBh
EHQqqcLwfMZOv2bLBwzZxP7WO7g7vcyZUd1aBlKZVap5OB5zEdTxfXnRoVY/73R7
ILOoOP6v6OLLiH8tqJmUe+pPR28iaakjAXiUjXpVWJs7Pj7E23Hr+5kGWrm03N0q
fDAY8py9j3kjyOEtd48KbWzx52wxNjwSE2AWxSHKrneX2KAibtxNLN8+K0iohfWJ
yP6zNsstXnH4WsE9C+xD/wz3PkFZ9m+s+d2GFXv17VgeDk/THJ8di2Yu8e2poRkU
vcxrVx/iYXdwIQYNfP2tFgc3ohbjKe7Er6NqZ0QHtFJdBFk4bogRN47OoWHyNv1Z
vlvOVzX2eTcV632JnoGe8Wx8UjhNJZRHQ+R/jog57AK8DcM6VeqMb5o57Ozd1m8/
by4XPYWhdXNB5Kdag6zW3r8KSe5BS+NoCn9BoRq/HR/QBt5RhTNaCbmY1DtYjWsh
U1029spsMSc0fvt50uV41Wx7FidliO+a5O1SSiuiiUggfzwdYV2usnZw14zsB+xz
0SShzblho6eXd5Sl/3OiitJDnM4aGJz8XYGqX+LDMslcOV01zbp1TrOS5Qjdlgk3
wb3N0WRH0b9d33kRczNAWykQTui+oEmq/rGQjcRzPBamNDgj9JF9FpcVZqY6tAIq
i2FdSIWYUgoPjYc1Wb0FDfuKOGoFFGMeV3cTn0spLTePBXVWhPQcezlaglcEE1CV
4nyVQDoLjUbeMwE5mziO6eREFpGzZC45RuKp9/S/WwfdQoOkFL9an9nI4t775GNv
jJxttcvgd9BEiK4J12E7P6kC7Wd58YLv/a4MTEVaFr9FwSjFz0fF2l6RRmC4HHCt
ekrKz4vlgaG6NFMo6LfrlC210CNwd8Vm4JKqP3VRpuhJFPqgK4tyrP+5mfQ8CT1p
9PZ/vKdDgKtAWzkQNyk+fxf7a+zEixIr9nGocbJE6pDTtpcOB+qGKRobSMBM1TtM
6ge3za7yuMJZuphZwR34MkAbKJFFQR+iSaHtCeiW3Z6KMBfu6StJzQqABKtkTBQO
ewXQs5j1X9PP9ErwkfzSW5322nmB8AvCK7KLyYhI/4vQkuxB00j7h9fTDS2n6F3Q
McDmfzLJ3SJIcViTx3OTdSD4IxF1EtM+KeUMH3VwWhx0oEao0UHJWFuM4xOebMz+
oBp4uDkvhGlXR4jBJs3g7+RVG6/Vp1bNKUeK6rCU+5LFonTvSxslgzIN0m6cYzxz
MGk9tpsfe8OgxzSel7Pmh8ASFO5rY/zJs0OMYPU6jKwoMH48l6aNLhz88f7+0T4n
eVWme/BBPOKQHqCYc+x/6G6rTwerSxXotdvhlqqJQBr7Vg8Ifp4LRwbpw1pH7azv
RjcTTu5+aVLtrhKTYRbYbuE9enVpNvqB31ibfEzYsFAcH4JJVz13XoEXepgJFDKO
AXwidGxqXQG/qLw/TqZ/tsLAq4YVhfE9i9Qm2FtZNU4VNjoWmALtzPYbMsTSm28B
IG9RWN/402MwV5BCo2ezblU873sNUmxIsQcJi9Zq/Y2ri0884wdmYdlAk/dGkajv
zhLLuKaeQmGGEpNURNATKAIU7ABUFKccLDH+3x4MlRAlpNay9FrHoT6Nl4aFpXDj
Pend5eOI+H3FR65Ket+3TUdRSjEzFLAyYvSydHZxvfqOmYqxtJ8kdUyXITmWzrGf
je5dlFVI/WOvkunCTs63jTtPI3ClMPsm35XPzls+HTZoieqL3WRjne4T916TO83+
GygGGh8MyqHLWpe6t4oe0FG67+NuI7cXlQT09kLzsbLiOIUdl3pnjVtMJg2yBy3w
tuIykpY4vsM+nUPSnkiuufRQmjWO8fD67szJqBnyA+RG2JaBcCjhoHYD5UDgElCY
ndvWUsVKYR4mcrGyAx44qS3UlbdkyrjMqCDUL9R18tZwzqnVdQetudadJEJQIGK/
InbnSepQyncBBJsHl4onzlOdoaiz23ZFnfnax7am2NMNGMFCT+++CsBXnmvfO3SF
NGuVvzaj9OdppgcfHH5hAR8TIyI49bIvUZG+Mx+ayWptXUhOGDUCSAYxUoroEBaN
Jdjc+pmObCTXNiCl9iuFRaDHjEGgDKoQ8wWCs/OCcm4+Q9iZ9eKO1iVmqojTgxse
riqcTah9XbPhQQIHVcztPo0ephjuJgdXJrLxEOa8JS9QW7z2L6DxKvQwpNaMicZO
VpDDH52awk+/io/pKWpXQgGUxubgOJiotohh+FlhRnYX8jk8ou1dZ1BjzCMc/lvJ
KgAq3BUT2GF9ScXYW1Jv4GIkXHdYeJrpqNUbkF6tx4YABjl7aJWWf7W1Vc/tsPG+
d8zuupJrmTVHpMrm+QUvmgl6RYdotbTv0dTy3DVzL5ZALckZissssYddp4QpMP96
uFbZIpfWQ4jXWhul6pdFR7L+2EiKVXn6Pqfr6caymwtCyILSJ/lbxMMGxDjbkU1L
h5KyWCngaKG/v5GJBRPvSpAjnOFXsBLodavRGoChvQwjq5sn/gKOPsE8KHfeuJH8
6MhKR/V0CyztehJ07yow4IPWSyVxuGihaAy/+FSmQiE8Lth4EJNN0vWXNRzcx1zl
0E2z7+I3hy+AzV6zo4QKAOfwLrR2ZD3cWtPKA5OVT4tIUSUxZ4CH35G9avNhEuw2
/P2Ku4Ycwcba3Q1vhk3YWsSTveMlx5h7OA2x6EMcs8Wca1m9H4fx5qkVRy1qn0Xw
zG0Kq0kkW1M0Rs8UT0Aj16No61MWHfxmxCWNWhbBQIJ+P2R/ohkRje9wSAnQr3wv
5sS1TlwAQRTBjhraSXpkh+8M/fqGJRYCZXj2Aywl8iC8L9FJ5ukRgF95Ukg47dQu
SZWxAuAJt+408K8IhBQbkKj3LwkvueqdEEtxpHHs/E+09B6mWsDNBlFqOgEOEqZG
idZ5nYoIfDwiU3Ej4o+29oMmKil/9jRx3hrgRm2guKSVBVJyCaozpfWvgurFkMks
E1qD5YMkH0q6G/0ikjrG3Kic2Fw07myLDiQzQxq5sDo49mOezxly2QxL+nXzr41h
GSPArP+KP55NR2MpEbCrWYT7ffpwdvP/H8DL5e/WNTYJjbDlaDOfJxc9p/nX4ILl
T3vcTFDS5HBSZrDZpXVJ/hc/1BqeMzeAiPlZGvL2ssEU4oealhEFZq8gSTKNwHkN
snU5BjFGikJJUf3Xd0Wm00Vme/CFKdwW+tDY74JVC8qMsik+qBX+KT+jwLhyTaOI
3o0mAiR7h0eJm6ondNn0WXGHBE5L2bpzKIw3+4qsD5sD8LKCE5cy23xrez2eC8Y7
14V4zPmJq6TQNTD0JwsaN2keRWCT7waVnkVn7wEhQAy/rYyP6K6r/47WqoZoBcl+
yC9v9gYRT95ouoG4MaveGrXuXCDkJKN0/JfGSoR4XOv49OZA9ZWjntfJEbmZZu+k
pV1sDDUIT7ThLGN0bgIxfJAP0EZjsDeBLhj2v/ZOICsnCXB7fGK9wcOGQw8N4JIW
zyvt/zGk1DTx66jCJAK0FdpizDbrZseDmHBKEkhg3d2FCGqe9FzLWdIrCgRSfKvg
1HB6jkfVtlVTAvYom9PDafzinVVahBRr5jmyzxpwjvBM0gz2z3DORzdT4bE27XKE
ZXJjA3320LpsizbLpxLGbLAhKxkmUEBZDh2VMmoUNclqtwwokSh21Xl/uCH4YUqi
gbndmHS+qjGnEsqXhZWU9rcy1RX0//bsVVxVD0E3dpMyb/bBsjH62EwK5z1MI0Jq
Fs5r78TiUJceX25s+dXJL7pSuWeAVDhD7jhMN/XItrU69LAwKrQx8eVeQNRvL97b
DXB2siFMZ2bKrjfYJnlQPTGZ7DiJHfjz1odqMb3w3KxpvwHiKrEnm7FYwoGOlG5z
YqN93JVaxLimmLog8VdEQqgW6Z3N7SMn8e91Z2AImUN1O5yDj+xfMYA6ONM1Nl7U
bN8l7WW7BeoA//PtiZ3oh6lbW8CteG46vsnTLjz5HSEmZ1DrBYJfYdcwH+dnPNgB
FjFFK0839O4S3IKuJeMHwlNm2JCKY6b7oQeyqHJYxr8CX0o1iGfh5pVGk0BwYKPn
U7Sf+13r6j7lD2XJ/BHhTpoX6Bx0J7If7UXuMLMVm+L36E4hwuHRtgRe6RQpgg5q
hBJ0GlJTBFybl8gPGd01B+kqVSj5MWRwsEY/4RGESoFngi67+ZvweJNqi3xLas0R
2U8q0txqRGIMnaMuBlcE85jjKvPmWYKjxrAPml0peWpUUDzs/2STpvkMwDjraxvC
jzaNmVZb9Ye7MfC8G6TPnRJyISgHPjyLlBB+ydBEKdiBM4Y3EgsXiOQjbemJX8QB
+KM6YoeCq0KIeo3oUj+CVNDji2f+0S25CNmfOUP6d49QnqsMcwrvr+bJOZfEEYt8
uDoH+2f4Oio3KuGjyRD82c4Exdolb5Z3NM8OVdjTIwzsmrWaWWevIqkuWlMpJwi5
4tS8f6TsvwOvT8NJ5WLcFTudceE5AQqpK/PoFJF1I95AW+h+KlOdXEmvcUv/titL
bQRNdVsRTl0mbVYUuWBRKbSe8cEne7P5Le9tT5an2VMwriEJLXZuy4e+sdzWxsrt
cLxSxZJmOxtYS0qzivzZdmadSU5boqL8xlBDVLsh6P41nZxFEtSa9/20eNeQ1V0j
+HxuIKrIrJTOOI8qOAYe5wnOcIBQY4hEVhPZtTg7jsztQeMKW9DX2wP2m89e0hKz
CLckpqnmDh0G/1RiBc5F8siZ6gDhnEysgHLJECXuFHB0kNtabtTqqEgLSo8uUoj3
2954mzNGbW5m/QBD/MawdYCBTtFXZeQjx9U84wO1UH0laMMleeBjhq0cOmAlwFzS
Oj+ETQvixYhkDYzqpdkqVZi7VQTR56jNlzRh4HFrd7fbysOfqygB/akOUfoADD2Z
AzsXCg7Lywuxiu/K10L++A==
`pragma protect end_protected
