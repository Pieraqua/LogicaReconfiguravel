`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
24ADmqn6lT6yHVXjsajdnnPQNEIi7Hp/Gj55iH6HTmnQGHSpiv444yBvCGrnGvlK
IcqwCg/FxQ1hvaNmCZRE22MOhEvnmijgNL7NHo9t/yIIpv8swaUYYsI9LZStQSVc
8G1ZrcOAbRkQN8617bgDV9eVbt7+jcz+eBLdylOV50ytkxsPFUG4tQlFqqpdsFZS
MfkPFVnBgjOnQ5iD6nV7cks/XENxjHeY/VcyKFLt5HTt+zIw/PMixCka6f0cSV8Y
wWkl3OEyr2R+jBLOgvBMULesC5lrUWRGg9o9PLqRnkwdfh0Gv1Rx/9jw9mdpmoiH
2+4tt5PcGP2g9qgYOYrX6QdU0fqjoyaRpBIIaBTrgNEIsMEZqnDolT3vFj+4p95b
jogBrWY0aPH+xFD+H9CNx80yNI+pT9pNIznXsWJNDW2EN5POC//mUR5YUdVy+2JJ
z9hfrA049USXjXhKFSeEx+tPlwKBi82zuuE4sGsWJ0K2HVI+OeMJehVkn2xsLs1q
hJfpFdjdMzVolOKUL+8Gylxue1fzJ1iYF18klYrzMMFomleg47iFvnE/WZUS7IJI
Fgbeh2TG+1WywGtQOBCVohz6yWEo2DijB4toJvWuvHiVeZTIRyj2ynuMvdrviFN4
JclPtT8XeygegmuaRwRxgdS3mthYmxtO0/w0QfKG/KhW0bv5PPONLv4qDzhunLxk
gPqaD/I7DPW+cqS4xNVLuvXXNBn0Odh/Nv495iArtLBuGArrLXK47kaf/pUkDxfj
OyR3zF0O23Sgto9GZIfh67l65N1f1E+tL3Qtp7p6d+SHECr85RVgt+hcum6H64DC
Kx9LY8gwsAI1FJBi8PMsgL08rZ67HXS6BmPblT7LMcC2WhKFEnnPGBVvwvEP/dJV
Peo8oo08MHHsOQOTfdg0RWINrb0IiedM9ON9MlAWEQ1tbX6q8dcygzB9py0xT/Jo
+9/heWWlg7e177eFL1zOlv8JQd7eb0ed4iPRXdRkCTLaa0nvMxLYrJLgioOyXLEr
/6tpniqsSi6aZorlWUV/s9zlTRVyOCeBF00XE3R2nxIUraHV3waBrgD2z8NhyUBo
5Q9WrkjI4nSIu1quktV/U2Dbn75+WlIdGtEZ2xzBaEyWLQxkbQRL2ZqvKGr0oTpR
x+MzpwPsq0k1oZL2KwOpABjI853DGxDJV7y9Lxwxqh5bLVNA2M7TuKZrBHkC9eE/
fvIgAkdD+p9q9EoY3YOJvpgQzEtM3acL+904a4ax2+TLRr5M5kS/mxbZ1m/3ae3W
dP7VJwRGguZwDc8j/iFUq/1j6vudOoCbid/hwrKX9t4Z2RTASsaQiG8xDXpOKdRj
rUWYMLTHVhvVB7zaTtceQvnt5BBo60G1ZDdZPZC5R4ykLNaa+qoaYTPAdI5Uxo8o
Fq9rCNdjCWlpNXAYJyE8KS1r4zsmU1imA62aUe0I8DqDGJROfGeCdp7JBvpU3JXg
Jpp8xQzsxh8O2O7tb8YYE8wwWg7WXskuvQJQif9HVm42ze0/Go+GSx7fraShbAG7
9wP0V5iEXVYxgtNSerucdL8/pRixVwdYt1PGp9SnQ4+Rla/6aRQt3NE3J6BHEKwG
eYgCpVbv8ZbZhCdUU5urRK1J3GKIJO8UTLL6JpUcE7NB0u/RFrT7Xl5VB9Je0/Po
F232YFys0UZOeYT0XosYcz1xCjUcGMHuXH57320wzYu91cYOwLQ6z4ZXj7HIGbVG
OaCngoD/bI0qSBE18eU4U4usAAnWuW/WYYlMO/FUlozeKffJxfhgofdNVh+7pNIR
6thbki/P6mFZgMD9uAEFDJuu14WwW9EzuULRGnYKkkKnmxkdjtGejH+i7YXnp89A
8PM80zl0YsnqYm3lumScE3Blducei8tTmgUjTEWypoTyF4MTLHefFjJbjAjpw8Oj
dq8yOptNRDoii5zjT+E1HbzeITzppbmSZSNWUwDFIHLAHxTUVaqub3AHPhnIVUnD
l7mI9CI3BmJF3KbSy/iEmpEYqPguO7FAi/nZosE1uLp6/acO5JFQ5jUXkeq1utk8
1uzObk5kV+LcKnu07M6w/bunueA7daQPb0jcd67xbu64cPgOwE6eCrZtb7B0dofy
6VNEIc7FRTWKwBgmYFEelTYhZnu3F27ICWVKCneQb8lOhUuwMgL0KBT+fqB6vf2x
ZFhsKwdjtcuWndkvOmY70XgvTymog8Qs3w5f27E0NYZ+NI1HnLkRcgFzDwDfIzxc
JXtG/4tb3b4r5TB8PITXAmqo95T7nJHUrH8vDW1JA7wxkhrNzM4c5pftmAB2Y4aK
oDJRvuGEDbKRsm66ptoreW0465mAQjuua+PzQMh8tZZXn1FDczABFIKnBw4g3/e6
II8gpeSwUQv/WczY5ke6V7qq4iSLGigcdQ58LVVaHgwvchA/RZjRlorWxGWYVHYS
NzBeVFTWPxoK2cAZLuWf1rSCRbUbqdJlSdCh3pE8hTwrmYyVSWx21t+sEb0c76DH
Fm9HM00IFZaUulPjCsRede9MMOBZ34ty+Chxq+s6C8lth7Plp2alWYLGLX0iCs2x
dphEHrJ4MBNMhy0E+wbyKoIl4C7++AN+euP1v3St+udUyDbGctcmt/hAd9MqlFwI
VRRx7sEHc5NZAiy+iB4aXnuvUI/oNrjGl5XeyjHnU8nuWfmJ5C3XBw5XktIs5oeG
X9Tn/6iOpOBs0OT5kp0dp7xkylUxD3D8aqrXK6NjBIlyDSHW+wKzqGjdvtTx+NPb
hDBrDJ3rMO8VyT8vBzwd6DeJU+VWHt29WJSXqHaYHpBH9n6VHhSG7E2tunU8L+zX
lwmRPYxO6iDi+WJnHDfDMiIOl9jj9Pa8JGCBaZ51DE3ladro9l25+ovzFTQfmvSz
iFZDQlkhATrQH/NP8YAqjNqf0iqBB2PHmeEb8zsSQoniB3bT7pUZWR+Wxz/9ys+5
L71BjvYFp9y3c1HvX1LyEA1dv+ZvLwE1Mr6eUgsVq8MyPPbB478gfu+FJSp2cP8v
BASk/PWMAmlQZWYzsWkSxkwUw4VHM/yTDriZKiFCnh0aJRF6m4z/KwJflsBLBHPc
cw/pnslHK6/yseNMXvIhUUxnYxXcOO63epETMjn+STvSU8wXfu2ZCkvPNGG+sLc4
fMJ0EvR3/qi+OVRO4mQ1XTRDGyAwNhXv2aoUKG5/Y3OAxHLIjDAPzi17ecOoyjH1
xbFK6PpCrvdutqjJ45wy96F1XpnBmsaRlE+/B077rd30Aa12tpY4upBPNmedPeCB
C4i0sDvtAn4XpAZkeWuzh1cZlpvCk/E+Bt5rBMZvhzfS2FXgvbc54r7XfKiFAJuh
XrjGn/OHoUP7KKFPwvGWACj0SAHUZ/dcGX/64JCN0hvhYDXwULdnKNRP6Lh1ZeEL
pSmN7HSxiZaiBqGmTWGto1VsNbSTuCjKs0G5x7LKv6eE9Ysjelbujzcb5O+sA4cA
NGoEr+GJ0J67qgQOEKkSHPP8Fqyg3tkRBdkNA62qrjxm8Fo+RbDcyEfQiTksgM9j
dvRrjFTO1/o2ZkbAfEZKkfStDx1Iw7Ve+SpKYBxW78/yIsM87TivboJ0NALuZXZE
X81VxfqCT+/z8u8XF/sV6ggEHW+QfIe1zBqE3ary8zBr052XeXI22KiU2pMc4+XE
cQbPVGeycvkhI3VqPFLTFdGTddppVfa4lWbpCgw0zqNp40Fm3ckrNoHnNEukrzBJ
nlsTDAYXqJGQEiRXeWLdUOSLdBz03hhx4lNHMc8pdOIcl7qb9WN1Sz68Xh+T7fvF
kw/Hxxiaz7EwMQn75ruIJNb1dMtgcINDCtXfsUhGwmXWab9dyDld1qqy+eJ68twu
M8wF+8iU0dkL/2ak2bJdmp1AT0jLad+u7p30YQFhgf4LPZH33eDkg3wKJBBZ1KfF
Iqdtkln1EEZvl28Vp2J3peJRMwHJ2izByreUlTVuhSFFWLPHizeNGhqRuBGBaDR7
9LKCmj4qdhXWFK7ByUhKVxg8S040Dv6Hn9chl5CrjUrRlgekk9/hmnVq2OgJFCDU
wHa4mjgW8/n+ZMW+gEM7JJY0hyXrknkc3aPa7gMIYlYb5V2EAl8tdk9HgAXp835M
7KO3sFWEMFymtDFx1wDXUxU7UOJc4hAQmlVKN6P2sHP3oVwtr7FFKWvvYDRLC4lL
x5601RuNBf/IR5afQDZxXeymcskJwhdATitVxbUBpBJ/IA7bpZ/K86YXTsfaVQ74
kzO3rwsrHbL41Wi5TksM6Ft6cSsAM3vL5C4dTdGj7VmdwAFwZh0aHBMuBXWw0/n9
GXunDN8qQGVv9vKbAPsdR6ZqDHlp7MmH39w4RCW9iAgb9AgpuuHwdOJieJ7LyNO7
VlFX7pm1xclCAOtiwUK8EZwitw8j2he0B3SpFBXwMViHvLZ4kj6cR+guLEfLHiNd
5T1SPoui+cz5TytRSdv94NfQu6j0fkNnUP/pTWe5VWMJA1JIbQm1R/ZQwYQoA6vf
cZD3pmnMxaRshuCUTzIER1M3HIEYMbeQccM67H4oDomUUEBtvctZkSy9HEDpfduC
k7WHy1anc/xLkhszrfp8Iyq54OOTPOAaNxTGtxZcrxlG1gm4mhZQjd8/DroATJIc
zvy9JI8NIwOYeCqdYotg8JseTVXB+gBprTRDfkGxQMMP41ORXVFvu0Ku6aRh6hSF
GP/OC65DBMBCg29juifvrgTcxSwuJFY1YojTqYt+5EFlteH8nOoUsu7y/7DiwrDT
lnAPKK98fFzsJFxfImMJexCrl/LK1dYKf/5qt2SgVG15olO9B/G6djQ/HI4NBUEu
TKdKyt+9jC8eSIavYN4x+wJ4mM/Tll/vNoVyJ0wIZ4ArMN4fPa4IZ474HoCj7x1r
PglVPdsB/sDZUDgc0un+DiLK2RSJA50/TOwlO5NX0g/LNF9shc+yIMs9HlPWWCTP
IBUpMYq/qkeJYxTYjJwSg/Bx67WeEoKduuObzi33uKe+DHV9zPJKZ8JN3fsEaQV3
vBwn4hFl3+6Ieu2G52YnLnJefOojhdAOnYvymadLjL8dTLVnwUY1Uv7c9Q+SdZb1
MR9Hkcyodh2kH2c05xWTbfDYRLByLKl3cB9BTFqGQuHKz2lxZbgHWu96jkOEe6ZZ
8/xAjVY6BmAS1GjbPaZJWwzjhhAdR/7KZ+efSrYtertSg4aVrLtRXrm1LDVuws/T
KRN9AFaxv48vKZGY4vM+TVsJ7ukMgbq+z3bQwESv0E5ZzbG986BEwXS0OdTiSiJA
yPqJrhWbVBogGqnnIalENNJAuV68W8uumwgMaTnRPyXtcbkX+CgUUI2+JCqncCRc
4mxrdUMETDGE2nImxJevwUFuExrbkegsRJr1DugV4Tl4mgj0Ead9Y+4DTbvQoN/9
7S2htnOSFpupmRegzi9b8n6A4G+g5xus/lWJyCSexDVLSp75U/5Ab5bpSx69qxbe
U4nlh7yp/fpa0WvtZJCqHkCxCt7ZRcCbMmaghU9M1RcFgiFZoHt/8BjxQf4u/H9O
Zky4C+SZOfh4Y5bQEEOzNKfChNUhPkQpU96nSmNc6tf8ZhdO5a8JO6ykYsLIz3Jn
l+xO6LHNdwwWY+ffLcpPlQ/u99Z4inuFzGbURhAxZyBD/xINLoGGduTls6NjEMH1
iyKWKjOP0JCG7I0ft/E27SeTLRK5Aonq4e7EFGWQgLoeJhpHpyKMK5e6qZmDeO6O
69kPHzEqRm0U3SzMzcCJEPGq6Ik1muFYbMuvX/K24C7JeK8tPVrZRZL2mtmBp3Bu
DEQuq3z7I8svW9vu+uKRi4wTtj/gAtN/zYPi2oteJMnDjvdU4dU3ZjZNeOFps6k9
7UqDED9vkCwgU7aY557hnGNIRqEI25oPFsv8s8rhw+5RyFCiPQSitMg9W1JhXzoG
fV4LId4gexlThvbbWsscFlngqNWqDpcKlYKRgLLmYeNLv/nYSCgGBstGLGETVqKx
pne4qjxPGJanLugOzxnpsStUeBQpYOkZDcwVs9JFipRX0/8tGc47f6fiwgj+jMK9
4jJb00Z6Z5YrXsmaCA6863re0kKira3D2AaWre89TmJT/73lrtGqtXms7Miuc6c0
OYR15tv6iBOanuaWhvNt5tZkK6S62vGkK4c8MEZ7CaMqaOXDUsL3yFZQJGRDuRdK
3abin1MVxzklAISu1/bJiIyO6DHAy7E+2bOisflxX6r3lLE/BsNrkllQtokpIkBR
0hSdpwlWkgawmDX+PVT1iWko8oyyQnhkCCaVW9DulijhDDIECvETP0XjAEkp8cIs
nGnIz3pzxqKRoC7fc0kJSS/v7VAVdNsQU3mWY4bUS0rM6eaW6XQp3NAIMliRW8fQ
CEiXWOX7XRiJi/RAeQZKEKAoKEPw95DuB/dsggiT67FzpsNYe8lcba35n0TlYAw3
NwibwJNDxHHHQOO8qWfn6mw8jrqIHxJNhrL9HfLp+aIL7fjXqBe1KdtvAG60WpbH
D7IToGx23pV5TPWZx6SCWx0cOPMA0sOIwgpZxL4mKbl2Ijx/AeWfOPLJ1pUcKBn5
pdpVrBRuYWvr99/izZOljXZlSRXOrVFXOs/e+FO++zmG1JpkID2MIR49u4SS2RV7
BIF9rmXhlTwPdJDo0/7qW1r3rbgP7RhnQjpyYhtA1HtIoKe8eR27881zkda8vuvd
XOyyylkmQGC0KDl1X/2XZKn+y43pNUPGxE/Obg3hITI=
`protect END_PROTECTED
